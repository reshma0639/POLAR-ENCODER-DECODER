`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: FWC IITH
// Engineer: Electronics engineer
// 
// Create Date: 30.12.2022 05:49:41
// Design Name: polar encoder
// Module Name: top_polar
// Project Name: polar encoder
// Target Devices: 
// Tool Versions: 
// Description: Perform polar encoder operation K=200,N=1024
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// This is the top module for polar encoder
//////////////////////////////////////////////////////////////////////////////////

module top_polar(
    input clk,empty,full,
    input rst,
    input  message,
   output reg result_s
    );
    reg [1023:0] result;

    wire [1023:0] inter_0;
    wire [1023:0] inter_1;
    wire [1023:0] inter_2;
    wire [1023:0] inter_3;
    wire [1023:0] inter_4;
    wire [1023:0] inter_5;
    wire [1023:0] inter_6;
    wire [1023:0] inter_7;
    wire [1023:0] inter_8;
    wire [1023:0] inter_9;
    wire [1023:0] inter_10;
    wire [1023:0] encoded_in;
    
    imps frozen(.smsg(message),.clk(clk),.reset(rst),.empty(empty),.full(full),.encoded(inter_0));
    assign inter_1[0] = inter_0[0]^inter_0[1];
    assign inter_1[1] = inter_0[1];
    assign inter_1[2] = inter_0[2]^inter_0[3];
    assign inter_1[3] = inter_0[3];
    assign inter_1[4] = inter_0[4]^inter_0[5];
    assign inter_1[5] = inter_0[5];
    assign inter_1[6] = inter_0[6]^inter_0[7];
    assign inter_1[7] = inter_0[7];
    assign inter_1[8] = inter_0[8]^inter_0[9];
    assign inter_1[9] = inter_0[9];
    assign inter_1[10] = inter_0[10]^inter_0[11];
    assign inter_1[11] = inter_0[11];
    assign inter_1[12] = inter_0[12]^inter_0[13];
    assign inter_1[13] = inter_0[13];
    assign inter_1[14] = inter_0[14]^inter_0[15];
    assign inter_1[15] = inter_0[15];
    assign inter_1[16] = inter_0[16]^inter_0[17];
    assign inter_1[17] = inter_0[17];
    assign inter_1[18] = inter_0[18]^inter_0[19];
    assign inter_1[19] = inter_0[19];
    assign inter_1[20] = inter_0[20]^inter_0[21];
    assign inter_1[21] = inter_0[21];
    assign inter_1[22] = inter_0[22]^inter_0[23];
    assign inter_1[23] = inter_0[23];
    assign inter_1[24] = inter_0[24]^inter_0[25];
    assign inter_1[25] = inter_0[25];
    assign inter_1[26] = inter_0[26]^inter_0[27];
    assign inter_1[27] = inter_0[27];
    assign inter_1[28] = inter_0[28]^inter_0[29];
    assign inter_1[29] = inter_0[29];
    assign inter_1[30] = inter_0[30]^inter_0[31];
    assign inter_1[31] = inter_0[31];
    assign inter_1[32] = inter_0[32]^inter_0[33];
    assign inter_1[33] = inter_0[33];
    assign inter_1[34] = inter_0[34]^inter_0[35];
    assign inter_1[35] = inter_0[35];
    assign inter_1[36] = inter_0[36]^inter_0[37];
    assign inter_1[37] = inter_0[37];
    assign inter_1[38] = inter_0[38]^inter_0[39];
    assign inter_1[39] = inter_0[39];
    assign inter_1[40] = inter_0[40]^inter_0[41];
    assign inter_1[41] = inter_0[41];
    assign inter_1[42] = inter_0[42]^inter_0[43];
    assign inter_1[43] = inter_0[43];
    assign inter_1[44] = inter_0[44]^inter_0[45];
    assign inter_1[45] = inter_0[45];
    assign inter_1[46] = inter_0[46]^inter_0[47];
    assign inter_1[47] = inter_0[47];
    assign inter_1[48] = inter_0[48]^inter_0[49];
    assign inter_1[49] = inter_0[49];
    assign inter_1[50] = inter_0[50]^inter_0[51];
    assign inter_1[51] = inter_0[51];
    assign inter_1[52] = inter_0[52]^inter_0[53];
    assign inter_1[53] = inter_0[53];
    assign inter_1[54] = inter_0[54]^inter_0[55];
    assign inter_1[55] = inter_0[55];
    assign inter_1[56] = inter_0[56]^inter_0[57];
    assign inter_1[57] = inter_0[57];
    assign inter_1[58] = inter_0[58]^inter_0[59];
    assign inter_1[59] = inter_0[59];
    assign inter_1[60] = inter_0[60]^inter_0[61];
    assign inter_1[61] = inter_0[61];
    assign inter_1[62] = inter_0[62]^inter_0[63];
    assign inter_1[63] = inter_0[63];
    assign inter_1[64] = inter_0[64]^inter_0[65];
    assign inter_1[65] = inter_0[65];
    assign inter_1[66] = inter_0[66]^inter_0[67];
    assign inter_1[67] = inter_0[67];
    assign inter_1[68] = inter_0[68]^inter_0[69];
    assign inter_1[69] = inter_0[69];
    assign inter_1[70] = inter_0[70]^inter_0[71];
    assign inter_1[71] = inter_0[71];
    assign inter_1[72] = inter_0[72]^inter_0[73];
    assign inter_1[73] = inter_0[73];
    assign inter_1[74] = inter_0[74]^inter_0[75];
    assign inter_1[75] = inter_0[75];
    assign inter_1[76] = inter_0[76]^inter_0[77];
    assign inter_1[77] = inter_0[77];
    assign inter_1[78] = inter_0[78]^inter_0[79];
    assign inter_1[79] = inter_0[79];
    assign inter_1[80] = inter_0[80]^inter_0[81];
    assign inter_1[81] = inter_0[81];
    assign inter_1[82] = inter_0[82]^inter_0[83];
    assign inter_1[83] = inter_0[83];
    assign inter_1[84] = inter_0[84]^inter_0[85];
    assign inter_1[85] = inter_0[85];
    assign inter_1[86] = inter_0[86]^inter_0[87];
    assign inter_1[87] = inter_0[87];
    assign inter_1[88] = inter_0[88]^inter_0[89];
    assign inter_1[89] = inter_0[89];
    assign inter_1[90] = inter_0[90]^inter_0[91];
    assign inter_1[91] = inter_0[91];
    assign inter_1[92] = inter_0[92]^inter_0[93];
    assign inter_1[93] = inter_0[93];
    assign inter_1[94] = inter_0[94]^inter_0[95];
    assign inter_1[95] = inter_0[95];
    assign inter_1[96] = inter_0[96]^inter_0[97];
    assign inter_1[97] = inter_0[97];
    assign inter_1[98] = inter_0[98]^inter_0[99];
    assign inter_1[99] = inter_0[99];
    assign inter_1[100] = inter_0[100]^inter_0[101];
    assign inter_1[101] = inter_0[101];
    assign inter_1[102] = inter_0[102]^inter_0[103];
    assign inter_1[103] = inter_0[103];
    assign inter_1[104] = inter_0[104]^inter_0[105];
    assign inter_1[105] = inter_0[105];
    assign inter_1[106] = inter_0[106]^inter_0[107];
    assign inter_1[107] = inter_0[107];
    assign inter_1[108] = inter_0[108]^inter_0[109];
    assign inter_1[109] = inter_0[109];
    assign inter_1[110] = inter_0[110]^inter_0[111];
    assign inter_1[111] = inter_0[111];
    assign inter_1[112] = inter_0[112]^inter_0[113];
    assign inter_1[113] = inter_0[113];
    assign inter_1[114] = inter_0[114]^inter_0[115];
    assign inter_1[115] = inter_0[115];
    assign inter_1[116] = inter_0[116]^inter_0[117];
    assign inter_1[117] = inter_0[117];
    assign inter_1[118] = inter_0[118]^inter_0[119];
    assign inter_1[119] = inter_0[119];
    assign inter_1[120] = inter_0[120]^inter_0[121];
    assign inter_1[121] = inter_0[121];
    assign inter_1[122] = inter_0[122]^inter_0[123];
    assign inter_1[123] = inter_0[123];
    assign inter_1[124] = inter_0[124]^inter_0[125];
    assign inter_1[125] = inter_0[125];
    assign inter_1[126] = inter_0[126]^inter_0[127];
    assign inter_1[127] = inter_0[127];
    assign inter_1[128] = inter_0[128]^inter_0[129];
    assign inter_1[129] = inter_0[129];
    assign inter_1[130] = inter_0[130]^inter_0[131];
    assign inter_1[131] = inter_0[131];
    assign inter_1[132] = inter_0[132]^inter_0[133];
    assign inter_1[133] = inter_0[133];
    assign inter_1[134] = inter_0[134]^inter_0[135];
    assign inter_1[135] = inter_0[135];
    assign inter_1[136] = inter_0[136]^inter_0[137];
    assign inter_1[137] = inter_0[137];
    assign inter_1[138] = inter_0[138]^inter_0[139];
    assign inter_1[139] = inter_0[139];
    assign inter_1[140] = inter_0[140]^inter_0[141];
    assign inter_1[141] = inter_0[141];
    assign inter_1[142] = inter_0[142]^inter_0[143];
    assign inter_1[143] = inter_0[143];
    assign inter_1[144] = inter_0[144]^inter_0[145];
    assign inter_1[145] = inter_0[145];
    assign inter_1[146] = inter_0[146]^inter_0[147];
    assign inter_1[147] = inter_0[147];
    assign inter_1[148] = inter_0[148]^inter_0[149];
    assign inter_1[149] = inter_0[149];
    assign inter_1[150] = inter_0[150]^inter_0[151];
    assign inter_1[151] = inter_0[151];
    assign inter_1[152] = inter_0[152]^inter_0[153];
    assign inter_1[153] = inter_0[153];
    assign inter_1[154] = inter_0[154]^inter_0[155];
    assign inter_1[155] = inter_0[155];
    assign inter_1[156] = inter_0[156]^inter_0[157];
    assign inter_1[157] = inter_0[157];
    assign inter_1[158] = inter_0[158]^inter_0[159];
    assign inter_1[159] = inter_0[159];
    assign inter_1[160] = inter_0[160]^inter_0[161];
    assign inter_1[161] = inter_0[161];
    assign inter_1[162] = inter_0[162]^inter_0[163];
    assign inter_1[163] = inter_0[163];
    assign inter_1[164] = inter_0[164]^inter_0[165];
    assign inter_1[165] = inter_0[165];
    assign inter_1[166] = inter_0[166]^inter_0[167];
    assign inter_1[167] = inter_0[167];
    assign inter_1[168] = inter_0[168]^inter_0[169];
    assign inter_1[169] = inter_0[169];
    assign inter_1[170] = inter_0[170]^inter_0[171];
    assign inter_1[171] = inter_0[171];
    assign inter_1[172] = inter_0[172]^inter_0[173];
    assign inter_1[173] = inter_0[173];
    assign inter_1[174] = inter_0[174]^inter_0[175];
    assign inter_1[175] = inter_0[175];
    assign inter_1[176] = inter_0[176]^inter_0[177];
    assign inter_1[177] = inter_0[177];
    assign inter_1[178] = inter_0[178]^inter_0[179];
    assign inter_1[179] = inter_0[179];
    assign inter_1[180] = inter_0[180]^inter_0[181];
    assign inter_1[181] = inter_0[181];
    assign inter_1[182] = inter_0[182]^inter_0[183];
    assign inter_1[183] = inter_0[183];
    assign inter_1[184] = inter_0[184]^inter_0[185];
    assign inter_1[185] = inter_0[185];
    assign inter_1[186] = inter_0[186]^inter_0[187];
    assign inter_1[187] = inter_0[187];
    assign inter_1[188] = inter_0[188]^inter_0[189];
    assign inter_1[189] = inter_0[189];
    assign inter_1[190] = inter_0[190]^inter_0[191];
    assign inter_1[191] = inter_0[191];
    assign inter_1[192] = inter_0[192]^inter_0[193];
    assign inter_1[193] = inter_0[193];
    assign inter_1[194] = inter_0[194]^inter_0[195];
    assign inter_1[195] = inter_0[195];
    assign inter_1[196] = inter_0[196]^inter_0[197];
    assign inter_1[197] = inter_0[197];
    assign inter_1[198] = inter_0[198]^inter_0[199];
    assign inter_1[199] = inter_0[199];
    assign inter_1[200] = inter_0[200]^inter_0[201];
    assign inter_1[201] = inter_0[201];
    assign inter_1[202] = inter_0[202]^inter_0[203];
    assign inter_1[203] = inter_0[203];
    assign inter_1[204] = inter_0[204]^inter_0[205];
    assign inter_1[205] = inter_0[205];
    assign inter_1[206] = inter_0[206]^inter_0[207];
    assign inter_1[207] = inter_0[207];
    assign inter_1[208] = inter_0[208]^inter_0[209];
    assign inter_1[209] = inter_0[209];
    assign inter_1[210] = inter_0[210]^inter_0[211];
    assign inter_1[211] = inter_0[211];
    assign inter_1[212] = inter_0[212]^inter_0[213];
    assign inter_1[213] = inter_0[213];
    assign inter_1[214] = inter_0[214]^inter_0[215];
    assign inter_1[215] = inter_0[215];
    assign inter_1[216] = inter_0[216]^inter_0[217];
    assign inter_1[217] = inter_0[217];
    assign inter_1[218] = inter_0[218]^inter_0[219];
    assign inter_1[219] = inter_0[219];
    assign inter_1[220] = inter_0[220]^inter_0[221];
    assign inter_1[221] = inter_0[221];
    assign inter_1[222] = inter_0[222]^inter_0[223];
    assign inter_1[223] = inter_0[223];
    assign inter_1[224] = inter_0[224]^inter_0[225];
    assign inter_1[225] = inter_0[225];
    assign inter_1[226] = inter_0[226]^inter_0[227];
    assign inter_1[227] = inter_0[227];
    assign inter_1[228] = inter_0[228]^inter_0[229];
    assign inter_1[229] = inter_0[229];
    assign inter_1[230] = inter_0[230]^inter_0[231];
    assign inter_1[231] = inter_0[231];
    assign inter_1[232] = inter_0[232]^inter_0[233];
    assign inter_1[233] = inter_0[233];
    assign inter_1[234] = inter_0[234]^inter_0[235];
    assign inter_1[235] = inter_0[235];
    assign inter_1[236] = inter_0[236]^inter_0[237];
    assign inter_1[237] = inter_0[237];
    assign inter_1[238] = inter_0[238]^inter_0[239];
    assign inter_1[239] = inter_0[239];
    assign inter_1[240] = inter_0[240]^inter_0[241];
    assign inter_1[241] = inter_0[241];
    assign inter_1[242] = inter_0[242]^inter_0[243];
    assign inter_1[243] = inter_0[243];
    assign inter_1[244] = inter_0[244]^inter_0[245];
    assign inter_1[245] = inter_0[245];
    assign inter_1[246] = inter_0[246]^inter_0[247];
    assign inter_1[247] = inter_0[247];
    assign inter_1[248] = inter_0[248]^inter_0[249];
    assign inter_1[249] = inter_0[249];
    assign inter_1[250] = inter_0[250]^inter_0[251];
    assign inter_1[251] = inter_0[251];
    assign inter_1[252] = inter_0[252]^inter_0[253];
    assign inter_1[253] = inter_0[253];
    assign inter_1[254] = inter_0[254]^inter_0[255];
    assign inter_1[255] = inter_0[255];
    assign inter_1[256] = inter_0[256]^inter_0[257];
    assign inter_1[257] = inter_0[257];
    assign inter_1[258] = inter_0[258]^inter_0[259];
    assign inter_1[259] = inter_0[259];
    assign inter_1[260] = inter_0[260]^inter_0[261];
    assign inter_1[261] = inter_0[261];
    assign inter_1[262] = inter_0[262]^inter_0[263];
    assign inter_1[263] = inter_0[263];
    assign inter_1[264] = inter_0[264]^inter_0[265];
    assign inter_1[265] = inter_0[265];
    assign inter_1[266] = inter_0[266]^inter_0[267];
    assign inter_1[267] = inter_0[267];
    assign inter_1[268] = inter_0[268]^inter_0[269];
    assign inter_1[269] = inter_0[269];
    assign inter_1[270] = inter_0[270]^inter_0[271];
    assign inter_1[271] = inter_0[271];
    assign inter_1[272] = inter_0[272]^inter_0[273];
    assign inter_1[273] = inter_0[273];
    assign inter_1[274] = inter_0[274]^inter_0[275];
    assign inter_1[275] = inter_0[275];
    assign inter_1[276] = inter_0[276]^inter_0[277];
    assign inter_1[277] = inter_0[277];
    assign inter_1[278] = inter_0[278]^inter_0[279];
    assign inter_1[279] = inter_0[279];
    assign inter_1[280] = inter_0[280]^inter_0[281];
    assign inter_1[281] = inter_0[281];
    assign inter_1[282] = inter_0[282]^inter_0[283];
    assign inter_1[283] = inter_0[283];
    assign inter_1[284] = inter_0[284]^inter_0[285];
    assign inter_1[285] = inter_0[285];
    assign inter_1[286] = inter_0[286]^inter_0[287];
    assign inter_1[287] = inter_0[287];
    assign inter_1[288] = inter_0[288]^inter_0[289];
    assign inter_1[289] = inter_0[289];
    assign inter_1[290] = inter_0[290]^inter_0[291];
    assign inter_1[291] = inter_0[291];
    assign inter_1[292] = inter_0[292]^inter_0[293];
    assign inter_1[293] = inter_0[293];
    assign inter_1[294] = inter_0[294]^inter_0[295];
    assign inter_1[295] = inter_0[295];
    assign inter_1[296] = inter_0[296]^inter_0[297];
    assign inter_1[297] = inter_0[297];
    assign inter_1[298] = inter_0[298]^inter_0[299];
    assign inter_1[299] = inter_0[299];
    assign inter_1[300] = inter_0[300]^inter_0[301];
    assign inter_1[301] = inter_0[301];
    assign inter_1[302] = inter_0[302]^inter_0[303];
    assign inter_1[303] = inter_0[303];
    assign inter_1[304] = inter_0[304]^inter_0[305];
    assign inter_1[305] = inter_0[305];
    assign inter_1[306] = inter_0[306]^inter_0[307];
    assign inter_1[307] = inter_0[307];
    assign inter_1[308] = inter_0[308]^inter_0[309];
    assign inter_1[309] = inter_0[309];
    assign inter_1[310] = inter_0[310]^inter_0[311];
    assign inter_1[311] = inter_0[311];
    assign inter_1[312] = inter_0[312]^inter_0[313];
    assign inter_1[313] = inter_0[313];
    assign inter_1[314] = inter_0[314]^inter_0[315];
    assign inter_1[315] = inter_0[315];
    assign inter_1[316] = inter_0[316]^inter_0[317];
    assign inter_1[317] = inter_0[317];
    assign inter_1[318] = inter_0[318]^inter_0[319];
    assign inter_1[319] = inter_0[319];
    assign inter_1[320] = inter_0[320]^inter_0[321];
    assign inter_1[321] = inter_0[321];
    assign inter_1[322] = inter_0[322]^inter_0[323];
    assign inter_1[323] = inter_0[323];
    assign inter_1[324] = inter_0[324]^inter_0[325];
    assign inter_1[325] = inter_0[325];
    assign inter_1[326] = inter_0[326]^inter_0[327];
    assign inter_1[327] = inter_0[327];
    assign inter_1[328] = inter_0[328]^inter_0[329];
    assign inter_1[329] = inter_0[329];
    assign inter_1[330] = inter_0[330]^inter_0[331];
    assign inter_1[331] = inter_0[331];
    assign inter_1[332] = inter_0[332]^inter_0[333];
    assign inter_1[333] = inter_0[333];
    assign inter_1[334] = inter_0[334]^inter_0[335];
    assign inter_1[335] = inter_0[335];
    assign inter_1[336] = inter_0[336]^inter_0[337];
    assign inter_1[337] = inter_0[337];
    assign inter_1[338] = inter_0[338]^inter_0[339];
    assign inter_1[339] = inter_0[339];
    assign inter_1[340] = inter_0[340]^inter_0[341];
    assign inter_1[341] = inter_0[341];
    assign inter_1[342] = inter_0[342]^inter_0[343];
    assign inter_1[343] = inter_0[343];
    assign inter_1[344] = inter_0[344]^inter_0[345];
    assign inter_1[345] = inter_0[345];
    assign inter_1[346] = inter_0[346]^inter_0[347];
    assign inter_1[347] = inter_0[347];
    assign inter_1[348] = inter_0[348]^inter_0[349];
    assign inter_1[349] = inter_0[349];
    assign inter_1[350] = inter_0[350]^inter_0[351];
    assign inter_1[351] = inter_0[351];
    assign inter_1[352] = inter_0[352]^inter_0[353];
    assign inter_1[353] = inter_0[353];
    assign inter_1[354] = inter_0[354]^inter_0[355];
    assign inter_1[355] = inter_0[355];
    assign inter_1[356] = inter_0[356]^inter_0[357];
    assign inter_1[357] = inter_0[357];
    assign inter_1[358] = inter_0[358]^inter_0[359];
    assign inter_1[359] = inter_0[359];
    assign inter_1[360] = inter_0[360]^inter_0[361];
    assign inter_1[361] = inter_0[361];
    assign inter_1[362] = inter_0[362]^inter_0[363];
    assign inter_1[363] = inter_0[363];
    assign inter_1[364] = inter_0[364]^inter_0[365];
    assign inter_1[365] = inter_0[365];
    assign inter_1[366] = inter_0[366]^inter_0[367];
    assign inter_1[367] = inter_0[367];
    assign inter_1[368] = inter_0[368]^inter_0[369];
    assign inter_1[369] = inter_0[369];
    assign inter_1[370] = inter_0[370]^inter_0[371];
    assign inter_1[371] = inter_0[371];
    assign inter_1[372] = inter_0[372]^inter_0[373];
    assign inter_1[373] = inter_0[373];
    assign inter_1[374] = inter_0[374]^inter_0[375];
    assign inter_1[375] = inter_0[375];
    assign inter_1[376] = inter_0[376]^inter_0[377];
    assign inter_1[377] = inter_0[377];
    assign inter_1[378] = inter_0[378]^inter_0[379];
    assign inter_1[379] = inter_0[379];
    assign inter_1[380] = inter_0[380]^inter_0[381];
    assign inter_1[381] = inter_0[381];
    assign inter_1[382] = inter_0[382]^inter_0[383];
    assign inter_1[383] = inter_0[383];
    assign inter_1[384] = inter_0[384]^inter_0[385];
    assign inter_1[385] = inter_0[385];
    assign inter_1[386] = inter_0[386]^inter_0[387];
    assign inter_1[387] = inter_0[387];
    assign inter_1[388] = inter_0[388]^inter_0[389];
    assign inter_1[389] = inter_0[389];
    assign inter_1[390] = inter_0[390]^inter_0[391];
    assign inter_1[391] = inter_0[391];
    assign inter_1[392] = inter_0[392]^inter_0[393];
    assign inter_1[393] = inter_0[393];
    assign inter_1[394] = inter_0[394]^inter_0[395];
    assign inter_1[395] = inter_0[395];
    assign inter_1[396] = inter_0[396]^inter_0[397];
    assign inter_1[397] = inter_0[397];
    assign inter_1[398] = inter_0[398]^inter_0[399];
    assign inter_1[399] = inter_0[399];
    assign inter_1[400] = inter_0[400]^inter_0[401];
    assign inter_1[401] = inter_0[401];
    assign inter_1[402] = inter_0[402]^inter_0[403];
    assign inter_1[403] = inter_0[403];
    assign inter_1[404] = inter_0[404]^inter_0[405];
    assign inter_1[405] = inter_0[405];
    assign inter_1[406] = inter_0[406]^inter_0[407];
    assign inter_1[407] = inter_0[407];
    assign inter_1[408] = inter_0[408]^inter_0[409];
    assign inter_1[409] = inter_0[409];
    assign inter_1[410] = inter_0[410]^inter_0[411];
    assign inter_1[411] = inter_0[411];
    assign inter_1[412] = inter_0[412]^inter_0[413];
    assign inter_1[413] = inter_0[413];
    assign inter_1[414] = inter_0[414]^inter_0[415];
    assign inter_1[415] = inter_0[415];
    assign inter_1[416] = inter_0[416]^inter_0[417];
    assign inter_1[417] = inter_0[417];
    assign inter_1[418] = inter_0[418]^inter_0[419];
    assign inter_1[419] = inter_0[419];
    assign inter_1[420] = inter_0[420]^inter_0[421];
    assign inter_1[421] = inter_0[421];
    assign inter_1[422] = inter_0[422]^inter_0[423];
    assign inter_1[423] = inter_0[423];
    assign inter_1[424] = inter_0[424]^inter_0[425];
    assign inter_1[425] = inter_0[425];
    assign inter_1[426] = inter_0[426]^inter_0[427];
    assign inter_1[427] = inter_0[427];
    assign inter_1[428] = inter_0[428]^inter_0[429];
    assign inter_1[429] = inter_0[429];
    assign inter_1[430] = inter_0[430]^inter_0[431];
    assign inter_1[431] = inter_0[431];
    assign inter_1[432] = inter_0[432]^inter_0[433];
    assign inter_1[433] = inter_0[433];
    assign inter_1[434] = inter_0[434]^inter_0[435];
    assign inter_1[435] = inter_0[435];
    assign inter_1[436] = inter_0[436]^inter_0[437];
    assign inter_1[437] = inter_0[437];
    assign inter_1[438] = inter_0[438]^inter_0[439];
    assign inter_1[439] = inter_0[439];
    assign inter_1[440] = inter_0[440]^inter_0[441];
    assign inter_1[441] = inter_0[441];
    assign inter_1[442] = inter_0[442]^inter_0[443];
    assign inter_1[443] = inter_0[443];
    assign inter_1[444] = inter_0[444]^inter_0[445];
    assign inter_1[445] = inter_0[445];
    assign inter_1[446] = inter_0[446]^inter_0[447];
    assign inter_1[447] = inter_0[447];
    assign inter_1[448] = inter_0[448]^inter_0[449];
    assign inter_1[449] = inter_0[449];
    assign inter_1[450] = inter_0[450]^inter_0[451];
    assign inter_1[451] = inter_0[451];
    assign inter_1[452] = inter_0[452]^inter_0[453];
    assign inter_1[453] = inter_0[453];
    assign inter_1[454] = inter_0[454]^inter_0[455];
    assign inter_1[455] = inter_0[455];
    assign inter_1[456] = inter_0[456]^inter_0[457];
    assign inter_1[457] = inter_0[457];
    assign inter_1[458] = inter_0[458]^inter_0[459];
    assign inter_1[459] = inter_0[459];
    assign inter_1[460] = inter_0[460]^inter_0[461];
    assign inter_1[461] = inter_0[461];
    assign inter_1[462] = inter_0[462]^inter_0[463];
    assign inter_1[463] = inter_0[463];
    assign inter_1[464] = inter_0[464]^inter_0[465];
    assign inter_1[465] = inter_0[465];
    assign inter_1[466] = inter_0[466]^inter_0[467];
    assign inter_1[467] = inter_0[467];
    assign inter_1[468] = inter_0[468]^inter_0[469];
    assign inter_1[469] = inter_0[469];
    assign inter_1[470] = inter_0[470]^inter_0[471];
    assign inter_1[471] = inter_0[471];
    assign inter_1[472] = inter_0[472]^inter_0[473];
    assign inter_1[473] = inter_0[473];
    assign inter_1[474] = inter_0[474]^inter_0[475];
    assign inter_1[475] = inter_0[475];
    assign inter_1[476] = inter_0[476]^inter_0[477];
    assign inter_1[477] = inter_0[477];
    assign inter_1[478] = inter_0[478]^inter_0[479];
    assign inter_1[479] = inter_0[479];
    assign inter_1[480] = inter_0[480]^inter_0[481];
    assign inter_1[481] = inter_0[481];
    assign inter_1[482] = inter_0[482]^inter_0[483];
    assign inter_1[483] = inter_0[483];
    assign inter_1[484] = inter_0[484]^inter_0[485];
    assign inter_1[485] = inter_0[485];
    assign inter_1[486] = inter_0[486]^inter_0[487];
    assign inter_1[487] = inter_0[487];
    assign inter_1[488] = inter_0[488]^inter_0[489];
    assign inter_1[489] = inter_0[489];
    assign inter_1[490] = inter_0[490]^inter_0[491];
    assign inter_1[491] = inter_0[491];
    assign inter_1[492] = inter_0[492]^inter_0[493];
    assign inter_1[493] = inter_0[493];
    assign inter_1[494] = inter_0[494]^inter_0[495];
    assign inter_1[495] = inter_0[495];
    assign inter_1[496] = inter_0[496]^inter_0[497];
    assign inter_1[497] = inter_0[497];
    assign inter_1[498] = inter_0[498]^inter_0[499];
    assign inter_1[499] = inter_0[499];
    assign inter_1[500] = inter_0[500]^inter_0[501];
    assign inter_1[501] = inter_0[501];
    assign inter_1[502] = inter_0[502]^inter_0[503];
    assign inter_1[503] = inter_0[503];
    assign inter_1[504] = inter_0[504]^inter_0[505];
    assign inter_1[505] = inter_0[505];
    assign inter_1[506] = inter_0[506]^inter_0[507];
    assign inter_1[507] = inter_0[507];
    assign inter_1[508] = inter_0[508]^inter_0[509];
    assign inter_1[509] = inter_0[509];
    assign inter_1[510] = inter_0[510]^inter_0[511];
    assign inter_1[511] = inter_0[511];
    assign inter_1[512] = inter_0[512]^inter_0[513];
    assign inter_1[513] = inter_0[513];
    assign inter_1[514] = inter_0[514]^inter_0[515];
    assign inter_1[515] = inter_0[515];
    assign inter_1[516] = inter_0[516]^inter_0[517];
    assign inter_1[517] = inter_0[517];
    assign inter_1[518] = inter_0[518]^inter_0[519];
    assign inter_1[519] = inter_0[519];
    assign inter_1[520] = inter_0[520]^inter_0[521];
    assign inter_1[521] = inter_0[521];
    assign inter_1[522] = inter_0[522]^inter_0[523];
    assign inter_1[523] = inter_0[523];
    assign inter_1[524] = inter_0[524]^inter_0[525];
    assign inter_1[525] = inter_0[525];
    assign inter_1[526] = inter_0[526]^inter_0[527];
    assign inter_1[527] = inter_0[527];
    assign inter_1[528] = inter_0[528]^inter_0[529];
    assign inter_1[529] = inter_0[529];
    assign inter_1[530] = inter_0[530]^inter_0[531];
    assign inter_1[531] = inter_0[531];
    assign inter_1[532] = inter_0[532]^inter_0[533];
    assign inter_1[533] = inter_0[533];
    assign inter_1[534] = inter_0[534]^inter_0[535];
    assign inter_1[535] = inter_0[535];
    assign inter_1[536] = inter_0[536]^inter_0[537];
    assign inter_1[537] = inter_0[537];
    assign inter_1[538] = inter_0[538]^inter_0[539];
    assign inter_1[539] = inter_0[539];
    assign inter_1[540] = inter_0[540]^inter_0[541];
    assign inter_1[541] = inter_0[541];
    assign inter_1[542] = inter_0[542]^inter_0[543];
    assign inter_1[543] = inter_0[543];
    assign inter_1[544] = inter_0[544]^inter_0[545];
    assign inter_1[545] = inter_0[545];
    assign inter_1[546] = inter_0[546]^inter_0[547];
    assign inter_1[547] = inter_0[547];
    assign inter_1[548] = inter_0[548]^inter_0[549];
    assign inter_1[549] = inter_0[549];
    assign inter_1[550] = inter_0[550]^inter_0[551];
    assign inter_1[551] = inter_0[551];
    assign inter_1[552] = inter_0[552]^inter_0[553];
    assign inter_1[553] = inter_0[553];
    assign inter_1[554] = inter_0[554]^inter_0[555];
    assign inter_1[555] = inter_0[555];
    assign inter_1[556] = inter_0[556]^inter_0[557];
    assign inter_1[557] = inter_0[557];
    assign inter_1[558] = inter_0[558]^inter_0[559];
    assign inter_1[559] = inter_0[559];
    assign inter_1[560] = inter_0[560]^inter_0[561];
    assign inter_1[561] = inter_0[561];
    assign inter_1[562] = inter_0[562]^inter_0[563];
    assign inter_1[563] = inter_0[563];
    assign inter_1[564] = inter_0[564]^inter_0[565];
    assign inter_1[565] = inter_0[565];
    assign inter_1[566] = inter_0[566]^inter_0[567];
    assign inter_1[567] = inter_0[567];
    assign inter_1[568] = inter_0[568]^inter_0[569];
    assign inter_1[569] = inter_0[569];
    assign inter_1[570] = inter_0[570]^inter_0[571];
    assign inter_1[571] = inter_0[571];
    assign inter_1[572] = inter_0[572]^inter_0[573];
    assign inter_1[573] = inter_0[573];
    assign inter_1[574] = inter_0[574]^inter_0[575];
    assign inter_1[575] = inter_0[575];
    assign inter_1[576] = inter_0[576]^inter_0[577];
    assign inter_1[577] = inter_0[577];
    assign inter_1[578] = inter_0[578]^inter_0[579];
    assign inter_1[579] = inter_0[579];
    assign inter_1[580] = inter_0[580]^inter_0[581];
    assign inter_1[581] = inter_0[581];
    assign inter_1[582] = inter_0[582]^inter_0[583];
    assign inter_1[583] = inter_0[583];
    assign inter_1[584] = inter_0[584]^inter_0[585];
    assign inter_1[585] = inter_0[585];
    assign inter_1[586] = inter_0[586]^inter_0[587];
    assign inter_1[587] = inter_0[587];
    assign inter_1[588] = inter_0[588]^inter_0[589];
    assign inter_1[589] = inter_0[589];
    assign inter_1[590] = inter_0[590]^inter_0[591];
    assign inter_1[591] = inter_0[591];
    assign inter_1[592] = inter_0[592]^inter_0[593];
    assign inter_1[593] = inter_0[593];
    assign inter_1[594] = inter_0[594]^inter_0[595];
    assign inter_1[595] = inter_0[595];
    assign inter_1[596] = inter_0[596]^inter_0[597];
    assign inter_1[597] = inter_0[597];
    assign inter_1[598] = inter_0[598]^inter_0[599];
    assign inter_1[599] = inter_0[599];
    assign inter_1[600] = inter_0[600]^inter_0[601];
    assign inter_1[601] = inter_0[601];
    assign inter_1[602] = inter_0[602]^inter_0[603];
    assign inter_1[603] = inter_0[603];
    assign inter_1[604] = inter_0[604]^inter_0[605];
    assign inter_1[605] = inter_0[605];
    assign inter_1[606] = inter_0[606]^inter_0[607];
    assign inter_1[607] = inter_0[607];
    assign inter_1[608] = inter_0[608]^inter_0[609];
    assign inter_1[609] = inter_0[609];
    assign inter_1[610] = inter_0[610]^inter_0[611];
    assign inter_1[611] = inter_0[611];
    assign inter_1[612] = inter_0[612]^inter_0[613];
    assign inter_1[613] = inter_0[613];
    assign inter_1[614] = inter_0[614]^inter_0[615];
    assign inter_1[615] = inter_0[615];
    assign inter_1[616] = inter_0[616]^inter_0[617];
    assign inter_1[617] = inter_0[617];
    assign inter_1[618] = inter_0[618]^inter_0[619];
    assign inter_1[619] = inter_0[619];
    assign inter_1[620] = inter_0[620]^inter_0[621];
    assign inter_1[621] = inter_0[621];
    assign inter_1[622] = inter_0[622]^inter_0[623];
    assign inter_1[623] = inter_0[623];
    assign inter_1[624] = inter_0[624]^inter_0[625];
    assign inter_1[625] = inter_0[625];
    assign inter_1[626] = inter_0[626]^inter_0[627];
    assign inter_1[627] = inter_0[627];
    assign inter_1[628] = inter_0[628]^inter_0[629];
    assign inter_1[629] = inter_0[629];
    assign inter_1[630] = inter_0[630]^inter_0[631];
    assign inter_1[631] = inter_0[631];
    assign inter_1[632] = inter_0[632]^inter_0[633];
    assign inter_1[633] = inter_0[633];
    assign inter_1[634] = inter_0[634]^inter_0[635];
    assign inter_1[635] = inter_0[635];
    assign inter_1[636] = inter_0[636]^inter_0[637];
    assign inter_1[637] = inter_0[637];
    assign inter_1[638] = inter_0[638]^inter_0[639];
    assign inter_1[639] = inter_0[639];
    assign inter_1[640] = inter_0[640]^inter_0[641];
    assign inter_1[641] = inter_0[641];
    assign inter_1[642] = inter_0[642]^inter_0[643];
    assign inter_1[643] = inter_0[643];
    assign inter_1[644] = inter_0[644]^inter_0[645];
    assign inter_1[645] = inter_0[645];
    assign inter_1[646] = inter_0[646]^inter_0[647];
    assign inter_1[647] = inter_0[647];
    assign inter_1[648] = inter_0[648]^inter_0[649];
    assign inter_1[649] = inter_0[649];
    assign inter_1[650] = inter_0[650]^inter_0[651];
    assign inter_1[651] = inter_0[651];
    assign inter_1[652] = inter_0[652]^inter_0[653];
    assign inter_1[653] = inter_0[653];
    assign inter_1[654] = inter_0[654]^inter_0[655];
    assign inter_1[655] = inter_0[655];
    assign inter_1[656] = inter_0[656]^inter_0[657];
    assign inter_1[657] = inter_0[657];
    assign inter_1[658] = inter_0[658]^inter_0[659];
    assign inter_1[659] = inter_0[659];
    assign inter_1[660] = inter_0[660]^inter_0[661];
    assign inter_1[661] = inter_0[661];
    assign inter_1[662] = inter_0[662]^inter_0[663];
    assign inter_1[663] = inter_0[663];
    assign inter_1[664] = inter_0[664]^inter_0[665];
    assign inter_1[665] = inter_0[665];
    assign inter_1[666] = inter_0[666]^inter_0[667];
    assign inter_1[667] = inter_0[667];
    assign inter_1[668] = inter_0[668]^inter_0[669];
    assign inter_1[669] = inter_0[669];
    assign inter_1[670] = inter_0[670]^inter_0[671];
    assign inter_1[671] = inter_0[671];
    assign inter_1[672] = inter_0[672]^inter_0[673];
    assign inter_1[673] = inter_0[673];
    assign inter_1[674] = inter_0[674]^inter_0[675];
    assign inter_1[675] = inter_0[675];
    assign inter_1[676] = inter_0[676]^inter_0[677];
    assign inter_1[677] = inter_0[677];
    assign inter_1[678] = inter_0[678]^inter_0[679];
    assign inter_1[679] = inter_0[679];
    assign inter_1[680] = inter_0[680]^inter_0[681];
    assign inter_1[681] = inter_0[681];
    assign inter_1[682] = inter_0[682]^inter_0[683];
    assign inter_1[683] = inter_0[683];
    assign inter_1[684] = inter_0[684]^inter_0[685];
    assign inter_1[685] = inter_0[685];
    assign inter_1[686] = inter_0[686]^inter_0[687];
    assign inter_1[687] = inter_0[687];
    assign inter_1[688] = inter_0[688]^inter_0[689];
    assign inter_1[689] = inter_0[689];
    assign inter_1[690] = inter_0[690]^inter_0[691];
    assign inter_1[691] = inter_0[691];
    assign inter_1[692] = inter_0[692]^inter_0[693];
    assign inter_1[693] = inter_0[693];
    assign inter_1[694] = inter_0[694]^inter_0[695];
    assign inter_1[695] = inter_0[695];
    assign inter_1[696] = inter_0[696]^inter_0[697];
    assign inter_1[697] = inter_0[697];
    assign inter_1[698] = inter_0[698]^inter_0[699];
    assign inter_1[699] = inter_0[699];
    assign inter_1[700] = inter_0[700]^inter_0[701];
    assign inter_1[701] = inter_0[701];
    assign inter_1[702] = inter_0[702]^inter_0[703];
    assign inter_1[703] = inter_0[703];
    assign inter_1[704] = inter_0[704]^inter_0[705];
    assign inter_1[705] = inter_0[705];
    assign inter_1[706] = inter_0[706]^inter_0[707];
    assign inter_1[707] = inter_0[707];
    assign inter_1[708] = inter_0[708]^inter_0[709];
    assign inter_1[709] = inter_0[709];
    assign inter_1[710] = inter_0[710]^inter_0[711];
    assign inter_1[711] = inter_0[711];
    assign inter_1[712] = inter_0[712]^inter_0[713];
    assign inter_1[713] = inter_0[713];
    assign inter_1[714] = inter_0[714]^inter_0[715];
    assign inter_1[715] = inter_0[715];
    assign inter_1[716] = inter_0[716]^inter_0[717];
    assign inter_1[717] = inter_0[717];
    assign inter_1[718] = inter_0[718]^inter_0[719];
    assign inter_1[719] = inter_0[719];
    assign inter_1[720] = inter_0[720]^inter_0[721];
    assign inter_1[721] = inter_0[721];
    assign inter_1[722] = inter_0[722]^inter_0[723];
    assign inter_1[723] = inter_0[723];
    assign inter_1[724] = inter_0[724]^inter_0[725];
    assign inter_1[725] = inter_0[725];
    assign inter_1[726] = inter_0[726]^inter_0[727];
    assign inter_1[727] = inter_0[727];
    assign inter_1[728] = inter_0[728]^inter_0[729];
    assign inter_1[729] = inter_0[729];
    assign inter_1[730] = inter_0[730]^inter_0[731];
    assign inter_1[731] = inter_0[731];
    assign inter_1[732] = inter_0[732]^inter_0[733];
    assign inter_1[733] = inter_0[733];
    assign inter_1[734] = inter_0[734]^inter_0[735];
    assign inter_1[735] = inter_0[735];
    assign inter_1[736] = inter_0[736]^inter_0[737];
    assign inter_1[737] = inter_0[737];
    assign inter_1[738] = inter_0[738]^inter_0[739];
    assign inter_1[739] = inter_0[739];
    assign inter_1[740] = inter_0[740]^inter_0[741];
    assign inter_1[741] = inter_0[741];
    assign inter_1[742] = inter_0[742]^inter_0[743];
    assign inter_1[743] = inter_0[743];
    assign inter_1[744] = inter_0[744]^inter_0[745];
    assign inter_1[745] = inter_0[745];
    assign inter_1[746] = inter_0[746]^inter_0[747];
    assign inter_1[747] = inter_0[747];
    assign inter_1[748] = inter_0[748]^inter_0[749];
    assign inter_1[749] = inter_0[749];
    assign inter_1[750] = inter_0[750]^inter_0[751];
    assign inter_1[751] = inter_0[751];
    assign inter_1[752] = inter_0[752]^inter_0[753];
    assign inter_1[753] = inter_0[753];
    assign inter_1[754] = inter_0[754]^inter_0[755];
    assign inter_1[755] = inter_0[755];
    assign inter_1[756] = inter_0[756]^inter_0[757];
    assign inter_1[757] = inter_0[757];
    assign inter_1[758] = inter_0[758]^inter_0[759];
    assign inter_1[759] = inter_0[759];
    assign inter_1[760] = inter_0[760]^inter_0[761];
    assign inter_1[761] = inter_0[761];
    assign inter_1[762] = inter_0[762]^inter_0[763];
    assign inter_1[763] = inter_0[763];
    assign inter_1[764] = inter_0[764]^inter_0[765];
    assign inter_1[765] = inter_0[765];
    assign inter_1[766] = inter_0[766]^inter_0[767];
    assign inter_1[767] = inter_0[767];
    assign inter_1[768] = inter_0[768]^inter_0[769];
    assign inter_1[769] = inter_0[769];
    assign inter_1[770] = inter_0[770]^inter_0[771];
    assign inter_1[771] = inter_0[771];
    assign inter_1[772] = inter_0[772]^inter_0[773];
    assign inter_1[773] = inter_0[773];
    assign inter_1[774] = inter_0[774]^inter_0[775];
    assign inter_1[775] = inter_0[775];
    assign inter_1[776] = inter_0[776]^inter_0[777];
    assign inter_1[777] = inter_0[777];
    assign inter_1[778] = inter_0[778]^inter_0[779];
    assign inter_1[779] = inter_0[779];
    assign inter_1[780] = inter_0[780]^inter_0[781];
    assign inter_1[781] = inter_0[781];
    assign inter_1[782] = inter_0[782]^inter_0[783];
    assign inter_1[783] = inter_0[783];
    assign inter_1[784] = inter_0[784]^inter_0[785];
    assign inter_1[785] = inter_0[785];
    assign inter_1[786] = inter_0[786]^inter_0[787];
    assign inter_1[787] = inter_0[787];
    assign inter_1[788] = inter_0[788]^inter_0[789];
    assign inter_1[789] = inter_0[789];
    assign inter_1[790] = inter_0[790]^inter_0[791];
    assign inter_1[791] = inter_0[791];
    assign inter_1[792] = inter_0[792]^inter_0[793];
    assign inter_1[793] = inter_0[793];
    assign inter_1[794] = inter_0[794]^inter_0[795];
    assign inter_1[795] = inter_0[795];
    assign inter_1[796] = inter_0[796]^inter_0[797];
    assign inter_1[797] = inter_0[797];
    assign inter_1[798] = inter_0[798]^inter_0[799];
    assign inter_1[799] = inter_0[799];
    assign inter_1[800] = inter_0[800]^inter_0[801];
    assign inter_1[801] = inter_0[801];
    assign inter_1[802] = inter_0[802]^inter_0[803];
    assign inter_1[803] = inter_0[803];
    assign inter_1[804] = inter_0[804]^inter_0[805];
    assign inter_1[805] = inter_0[805];
    assign inter_1[806] = inter_0[806]^inter_0[807];
    assign inter_1[807] = inter_0[807];
    assign inter_1[808] = inter_0[808]^inter_0[809];
    assign inter_1[809] = inter_0[809];
    assign inter_1[810] = inter_0[810]^inter_0[811];
    assign inter_1[811] = inter_0[811];
    assign inter_1[812] = inter_0[812]^inter_0[813];
    assign inter_1[813] = inter_0[813];
    assign inter_1[814] = inter_0[814]^inter_0[815];
    assign inter_1[815] = inter_0[815];
    assign inter_1[816] = inter_0[816]^inter_0[817];
    assign inter_1[817] = inter_0[817];
    assign inter_1[818] = inter_0[818]^inter_0[819];
    assign inter_1[819] = inter_0[819];
    assign inter_1[820] = inter_0[820]^inter_0[821];
    assign inter_1[821] = inter_0[821];
    assign inter_1[822] = inter_0[822]^inter_0[823];
    assign inter_1[823] = inter_0[823];
    assign inter_1[824] = inter_0[824]^inter_0[825];
    assign inter_1[825] = inter_0[825];
    assign inter_1[826] = inter_0[826]^inter_0[827];
    assign inter_1[827] = inter_0[827];
    assign inter_1[828] = inter_0[828]^inter_0[829];
    assign inter_1[829] = inter_0[829];
    assign inter_1[830] = inter_0[830]^inter_0[831];
    assign inter_1[831] = inter_0[831];
    assign inter_1[832] = inter_0[832]^inter_0[833];
    assign inter_1[833] = inter_0[833];
    assign inter_1[834] = inter_0[834]^inter_0[835];
    assign inter_1[835] = inter_0[835];
    assign inter_1[836] = inter_0[836]^inter_0[837];
    assign inter_1[837] = inter_0[837];
    assign inter_1[838] = inter_0[838]^inter_0[839];
    assign inter_1[839] = inter_0[839];
    assign inter_1[840] = inter_0[840]^inter_0[841];
    assign inter_1[841] = inter_0[841];
    assign inter_1[842] = inter_0[842]^inter_0[843];
    assign inter_1[843] = inter_0[843];
    assign inter_1[844] = inter_0[844]^inter_0[845];
    assign inter_1[845] = inter_0[845];
    assign inter_1[846] = inter_0[846]^inter_0[847];
    assign inter_1[847] = inter_0[847];
    assign inter_1[848] = inter_0[848]^inter_0[849];
    assign inter_1[849] = inter_0[849];
    assign inter_1[850] = inter_0[850]^inter_0[851];
    assign inter_1[851] = inter_0[851];
    assign inter_1[852] = inter_0[852]^inter_0[853];
    assign inter_1[853] = inter_0[853];
    assign inter_1[854] = inter_0[854]^inter_0[855];
    assign inter_1[855] = inter_0[855];
    assign inter_1[856] = inter_0[856]^inter_0[857];
    assign inter_1[857] = inter_0[857];
    assign inter_1[858] = inter_0[858]^inter_0[859];
    assign inter_1[859] = inter_0[859];
    assign inter_1[860] = inter_0[860]^inter_0[861];
    assign inter_1[861] = inter_0[861];
    assign inter_1[862] = inter_0[862]^inter_0[863];
    assign inter_1[863] = inter_0[863];
    assign inter_1[864] = inter_0[864]^inter_0[865];
    assign inter_1[865] = inter_0[865];
    assign inter_1[866] = inter_0[866]^inter_0[867];
    assign inter_1[867] = inter_0[867];
    assign inter_1[868] = inter_0[868]^inter_0[869];
    assign inter_1[869] = inter_0[869];
    assign inter_1[870] = inter_0[870]^inter_0[871];
    assign inter_1[871] = inter_0[871];
    assign inter_1[872] = inter_0[872]^inter_0[873];
    assign inter_1[873] = inter_0[873];
    assign inter_1[874] = inter_0[874]^inter_0[875];
    assign inter_1[875] = inter_0[875];
    assign inter_1[876] = inter_0[876]^inter_0[877];
    assign inter_1[877] = inter_0[877];
    assign inter_1[878] = inter_0[878]^inter_0[879];
    assign inter_1[879] = inter_0[879];
    assign inter_1[880] = inter_0[880]^inter_0[881];
    assign inter_1[881] = inter_0[881];
    assign inter_1[882] = inter_0[882]^inter_0[883];
    assign inter_1[883] = inter_0[883];
    assign inter_1[884] = inter_0[884]^inter_0[885];
    assign inter_1[885] = inter_0[885];
    assign inter_1[886] = inter_0[886]^inter_0[887];
    assign inter_1[887] = inter_0[887];
    assign inter_1[888] = inter_0[888]^inter_0[889];
    assign inter_1[889] = inter_0[889];
    assign inter_1[890] = inter_0[890]^inter_0[891];
    assign inter_1[891] = inter_0[891];
    assign inter_1[892] = inter_0[892]^inter_0[893];
    assign inter_1[893] = inter_0[893];
    assign inter_1[894] = inter_0[894]^inter_0[895];
    assign inter_1[895] = inter_0[895];
    assign inter_1[896] = inter_0[896]^inter_0[897];
    assign inter_1[897] = inter_0[897];
    assign inter_1[898] = inter_0[898]^inter_0[899];
    assign inter_1[899] = inter_0[899];
    assign inter_1[900] = inter_0[900]^inter_0[901];
    assign inter_1[901] = inter_0[901];
    assign inter_1[902] = inter_0[902]^inter_0[903];
    assign inter_1[903] = inter_0[903];
    assign inter_1[904] = inter_0[904]^inter_0[905];
    assign inter_1[905] = inter_0[905];
    assign inter_1[906] = inter_0[906]^inter_0[907];
    assign inter_1[907] = inter_0[907];
    assign inter_1[908] = inter_0[908]^inter_0[909];
    assign inter_1[909] = inter_0[909];
    assign inter_1[910] = inter_0[910]^inter_0[911];
    assign inter_1[911] = inter_0[911];
    assign inter_1[912] = inter_0[912]^inter_0[913];
    assign inter_1[913] = inter_0[913];
    assign inter_1[914] = inter_0[914]^inter_0[915];
    assign inter_1[915] = inter_0[915];
    assign inter_1[916] = inter_0[916]^inter_0[917];
    assign inter_1[917] = inter_0[917];
    assign inter_1[918] = inter_0[918]^inter_0[919];
    assign inter_1[919] = inter_0[919];
    assign inter_1[920] = inter_0[920]^inter_0[921];
    assign inter_1[921] = inter_0[921];
    assign inter_1[922] = inter_0[922]^inter_0[923];
    assign inter_1[923] = inter_0[923];
    assign inter_1[924] = inter_0[924]^inter_0[925];
    assign inter_1[925] = inter_0[925];
    assign inter_1[926] = inter_0[926]^inter_0[927];
    assign inter_1[927] = inter_0[927];
    assign inter_1[928] = inter_0[928]^inter_0[929];
    assign inter_1[929] = inter_0[929];
    assign inter_1[930] = inter_0[930]^inter_0[931];
    assign inter_1[931] = inter_0[931];
    assign inter_1[932] = inter_0[932]^inter_0[933];
    assign inter_1[933] = inter_0[933];
    assign inter_1[934] = inter_0[934]^inter_0[935];
    assign inter_1[935] = inter_0[935];
    assign inter_1[936] = inter_0[936]^inter_0[937];
    assign inter_1[937] = inter_0[937];
    assign inter_1[938] = inter_0[938]^inter_0[939];
    assign inter_1[939] = inter_0[939];
    assign inter_1[940] = inter_0[940]^inter_0[941];
    assign inter_1[941] = inter_0[941];
    assign inter_1[942] = inter_0[942]^inter_0[943];
    assign inter_1[943] = inter_0[943];
    assign inter_1[944] = inter_0[944]^inter_0[945];
    assign inter_1[945] = inter_0[945];
    assign inter_1[946] = inter_0[946]^inter_0[947];
    assign inter_1[947] = inter_0[947];
    assign inter_1[948] = inter_0[948]^inter_0[949];
    assign inter_1[949] = inter_0[949];
    assign inter_1[950] = inter_0[950]^inter_0[951];
    assign inter_1[951] = inter_0[951];
    assign inter_1[952] = inter_0[952]^inter_0[953];
    assign inter_1[953] = inter_0[953];
    assign inter_1[954] = inter_0[954]^inter_0[955];
    assign inter_1[955] = inter_0[955];
    assign inter_1[956] = inter_0[956]^inter_0[957];
    assign inter_1[957] = inter_0[957];
    assign inter_1[958] = inter_0[958]^inter_0[959];
    assign inter_1[959] = inter_0[959];
    assign inter_1[960] = inter_0[960]^inter_0[961];
    assign inter_1[961] = inter_0[961];
    assign inter_1[962] = inter_0[962]^inter_0[963];
    assign inter_1[963] = inter_0[963];
    assign inter_1[964] = inter_0[964]^inter_0[965];
    assign inter_1[965] = inter_0[965];
    assign inter_1[966] = inter_0[966]^inter_0[967];
    assign inter_1[967] = inter_0[967];
    assign inter_1[968] = inter_0[968]^inter_0[969];
    assign inter_1[969] = inter_0[969];
    assign inter_1[970] = inter_0[970]^inter_0[971];
    assign inter_1[971] = inter_0[971];
    assign inter_1[972] = inter_0[972]^inter_0[973];
    assign inter_1[973] = inter_0[973];
    assign inter_1[974] = inter_0[974]^inter_0[975];
    assign inter_1[975] = inter_0[975];
    assign inter_1[976] = inter_0[976]^inter_0[977];
    assign inter_1[977] = inter_0[977];
    assign inter_1[978] = inter_0[978]^inter_0[979];
    assign inter_1[979] = inter_0[979];
    assign inter_1[980] = inter_0[980]^inter_0[981];
    assign inter_1[981] = inter_0[981];
    assign inter_1[982] = inter_0[982]^inter_0[983];
    assign inter_1[983] = inter_0[983];
    assign inter_1[984] = inter_0[984]^inter_0[985];
    assign inter_1[985] = inter_0[985];
    assign inter_1[986] = inter_0[986]^inter_0[987];
    assign inter_1[987] = inter_0[987];
    assign inter_1[988] = inter_0[988]^inter_0[989];
    assign inter_1[989] = inter_0[989];
    assign inter_1[990] = inter_0[990]^inter_0[991];
    assign inter_1[991] = inter_0[991];
    assign inter_1[992] = inter_0[992]^inter_0[993];
    assign inter_1[993] = inter_0[993];
    assign inter_1[994] = inter_0[994]^inter_0[995];
    assign inter_1[995] = inter_0[995];
    assign inter_1[996] = inter_0[996]^inter_0[997];
    assign inter_1[997] = inter_0[997];
    assign inter_1[998] = inter_0[998]^inter_0[999];
    assign inter_1[999] = inter_0[999];
    assign inter_1[1000] = inter_0[1000]^inter_0[1001];
    assign inter_1[1001] = inter_0[1001];
    assign inter_1[1002] = inter_0[1002]^inter_0[1003];
    assign inter_1[1003] = inter_0[1003];
    assign inter_1[1004] = inter_0[1004]^inter_0[1005];
    assign inter_1[1005] = inter_0[1005];
    assign inter_1[1006] = inter_0[1006]^inter_0[1007];
    assign inter_1[1007] = inter_0[1007];
    assign inter_1[1008] = inter_0[1008]^inter_0[1009];
    assign inter_1[1009] = inter_0[1009];
    assign inter_1[1010] = inter_0[1010]^inter_0[1011];
    assign inter_1[1011] = inter_0[1011];
    assign inter_1[1012] = inter_0[1012]^inter_0[1013];
    assign inter_1[1013] = inter_0[1013];
    assign inter_1[1014] = inter_0[1014]^inter_0[1015];
    assign inter_1[1015] = inter_0[1015];
    assign inter_1[1016] = inter_0[1016]^inter_0[1017];
    assign inter_1[1017] = inter_0[1017];
    assign inter_1[1018] = inter_0[1018]^inter_0[1019];
    assign inter_1[1019] = inter_0[1019];
    assign inter_1[1020] = inter_0[1020]^inter_0[1021];
    assign inter_1[1021] = inter_0[1021];
    assign inter_1[1022] = inter_0[1022]^inter_0[1023];
    assign inter_1[1023] = inter_0[1023];
    /***************************/
    assign inter_2[0] = inter_1[0]^inter_1[2];
    assign inter_2[1] = inter_1[1]^inter_1[3];
    assign inter_2[2] = inter_1[2];
    assign inter_2[3] = inter_1[3];
    assign inter_2[4] = inter_1[4]^inter_1[6];
    assign inter_2[5] = inter_1[5]^inter_1[7];
    assign inter_2[6] = inter_1[6];
    assign inter_2[7] = inter_1[7];
    assign inter_2[8] = inter_1[8]^inter_1[10];
    assign inter_2[9] = inter_1[9]^inter_1[11];
    assign inter_2[10] = inter_1[10];
    assign inter_2[11] = inter_1[11];
    assign inter_2[12] = inter_1[12]^inter_1[14];
    assign inter_2[13] = inter_1[13]^inter_1[15];
    assign inter_2[14] = inter_1[14];
    assign inter_2[15] = inter_1[15];
    assign inter_2[16] = inter_1[16]^inter_1[18];
    assign inter_2[17] = inter_1[17]^inter_1[19];
    assign inter_2[18] = inter_1[18];
    assign inter_2[19] = inter_1[19];
    assign inter_2[20] = inter_1[20]^inter_1[22];
    assign inter_2[21] = inter_1[21]^inter_1[23];
    assign inter_2[22] = inter_1[22];
    assign inter_2[23] = inter_1[23];
    assign inter_2[24] = inter_1[24]^inter_1[26];
    assign inter_2[25] = inter_1[25]^inter_1[27];
    assign inter_2[26] = inter_1[26];
    assign inter_2[27] = inter_1[27];
    assign inter_2[28] = inter_1[28]^inter_1[30];
    assign inter_2[29] = inter_1[29]^inter_1[31];
    assign inter_2[30] = inter_1[30];
    assign inter_2[31] = inter_1[31];
    assign inter_2[32] = inter_1[32]^inter_1[34];
    assign inter_2[33] = inter_1[33]^inter_1[35];
    assign inter_2[34] = inter_1[34];
    assign inter_2[35] = inter_1[35];
    assign inter_2[36] = inter_1[36]^inter_1[38];
    assign inter_2[37] = inter_1[37]^inter_1[39];
    assign inter_2[38] = inter_1[38];
    assign inter_2[39] = inter_1[39];
    assign inter_2[40] = inter_1[40]^inter_1[42];
    assign inter_2[41] = inter_1[41]^inter_1[43];
    assign inter_2[42] = inter_1[42];
    assign inter_2[43] = inter_1[43];
    assign inter_2[44] = inter_1[44]^inter_1[46];
    assign inter_2[45] = inter_1[45]^inter_1[47];
    assign inter_2[46] = inter_1[46];
    assign inter_2[47] = inter_1[47];
    assign inter_2[48] = inter_1[48]^inter_1[50];
    assign inter_2[49] = inter_1[49]^inter_1[51];
    assign inter_2[50] = inter_1[50];
    assign inter_2[51] = inter_1[51];
    assign inter_2[52] = inter_1[52]^inter_1[54];
    assign inter_2[53] = inter_1[53]^inter_1[55];
    assign inter_2[54] = inter_1[54];
    assign inter_2[55] = inter_1[55];
    assign inter_2[56] = inter_1[56]^inter_1[58];
    assign inter_2[57] = inter_1[57]^inter_1[59];
    assign inter_2[58] = inter_1[58];
    assign inter_2[59] = inter_1[59];
    assign inter_2[60] = inter_1[60]^inter_1[62];
    assign inter_2[61] = inter_1[61]^inter_1[63];
    assign inter_2[62] = inter_1[62];
    assign inter_2[63] = inter_1[63];
    assign inter_2[64] = inter_1[64]^inter_1[66];
    assign inter_2[65] = inter_1[65]^inter_1[67];
    assign inter_2[66] = inter_1[66];
    assign inter_2[67] = inter_1[67];
    assign inter_2[68] = inter_1[68]^inter_1[70];
    assign inter_2[69] = inter_1[69]^inter_1[71];
    assign inter_2[70] = inter_1[70];
    assign inter_2[71] = inter_1[71];
    assign inter_2[72] = inter_1[72]^inter_1[74];
    assign inter_2[73] = inter_1[73]^inter_1[75];
    assign inter_2[74] = inter_1[74];
    assign inter_2[75] = inter_1[75];
    assign inter_2[76] = inter_1[76]^inter_1[78];
    assign inter_2[77] = inter_1[77]^inter_1[79];
    assign inter_2[78] = inter_1[78];
    assign inter_2[79] = inter_1[79];
    assign inter_2[80] = inter_1[80]^inter_1[82];
    assign inter_2[81] = inter_1[81]^inter_1[83];
    assign inter_2[82] = inter_1[82];
    assign inter_2[83] = inter_1[83];
    assign inter_2[84] = inter_1[84]^inter_1[86];
    assign inter_2[85] = inter_1[85]^inter_1[87];
    assign inter_2[86] = inter_1[86];
    assign inter_2[87] = inter_1[87];
    assign inter_2[88] = inter_1[88]^inter_1[90];
    assign inter_2[89] = inter_1[89]^inter_1[91];
    assign inter_2[90] = inter_1[90];
    assign inter_2[91] = inter_1[91];
    assign inter_2[92] = inter_1[92]^inter_1[94];
    assign inter_2[93] = inter_1[93]^inter_1[95];
    assign inter_2[94] = inter_1[94];
    assign inter_2[95] = inter_1[95];
    assign inter_2[96] = inter_1[96]^inter_1[98];
    assign inter_2[97] = inter_1[97]^inter_1[99];
    assign inter_2[98] = inter_1[98];
    assign inter_2[99] = inter_1[99];
    assign inter_2[100] = inter_1[100]^inter_1[102];
    assign inter_2[101] = inter_1[101]^inter_1[103];
    assign inter_2[102] = inter_1[102];
    assign inter_2[103] = inter_1[103];
    assign inter_2[104] = inter_1[104]^inter_1[106];
    assign inter_2[105] = inter_1[105]^inter_1[107];
    assign inter_2[106] = inter_1[106];
    assign inter_2[107] = inter_1[107];
    assign inter_2[108] = inter_1[108]^inter_1[110];
    assign inter_2[109] = inter_1[109]^inter_1[111];
    assign inter_2[110] = inter_1[110];
    assign inter_2[111] = inter_1[111];
    assign inter_2[112] = inter_1[112]^inter_1[114];
    assign inter_2[113] = inter_1[113]^inter_1[115];
    assign inter_2[114] = inter_1[114];
    assign inter_2[115] = inter_1[115];
    assign inter_2[116] = inter_1[116]^inter_1[118];
    assign inter_2[117] = inter_1[117]^inter_1[119];
    assign inter_2[118] = inter_1[118];
    assign inter_2[119] = inter_1[119];
    assign inter_2[120] = inter_1[120]^inter_1[122];
    assign inter_2[121] = inter_1[121]^inter_1[123];
    assign inter_2[122] = inter_1[122];
    assign inter_2[123] = inter_1[123];
    assign inter_2[124] = inter_1[124]^inter_1[126];
    assign inter_2[125] = inter_1[125]^inter_1[127];
    assign inter_2[126] = inter_1[126];
    assign inter_2[127] = inter_1[127];
    assign inter_2[128] = inter_1[128]^inter_1[130];
    assign inter_2[129] = inter_1[129]^inter_1[131];
    assign inter_2[130] = inter_1[130];
    assign inter_2[131] = inter_1[131];
    assign inter_2[132] = inter_1[132]^inter_1[134];
    assign inter_2[133] = inter_1[133]^inter_1[135];
    assign inter_2[134] = inter_1[134];
    assign inter_2[135] = inter_1[135];
    assign inter_2[136] = inter_1[136]^inter_1[138];
    assign inter_2[137] = inter_1[137]^inter_1[139];
    assign inter_2[138] = inter_1[138];
    assign inter_2[139] = inter_1[139];
    assign inter_2[140] = inter_1[140]^inter_1[142];
    assign inter_2[141] = inter_1[141]^inter_1[143];
    assign inter_2[142] = inter_1[142];
    assign inter_2[143] = inter_1[143];
    assign inter_2[144] = inter_1[144]^inter_1[146];
    assign inter_2[145] = inter_1[145]^inter_1[147];
    assign inter_2[146] = inter_1[146];
    assign inter_2[147] = inter_1[147];
    assign inter_2[148] = inter_1[148]^inter_1[150];
    assign inter_2[149] = inter_1[149]^inter_1[151];
    assign inter_2[150] = inter_1[150];
    assign inter_2[151] = inter_1[151];
    assign inter_2[152] = inter_1[152]^inter_1[154];
    assign inter_2[153] = inter_1[153]^inter_1[155];
    assign inter_2[154] = inter_1[154];
    assign inter_2[155] = inter_1[155];
    assign inter_2[156] = inter_1[156]^inter_1[158];
    assign inter_2[157] = inter_1[157]^inter_1[159];
    assign inter_2[158] = inter_1[158];
    assign inter_2[159] = inter_1[159];
    assign inter_2[160] = inter_1[160]^inter_1[162];
    assign inter_2[161] = inter_1[161]^inter_1[163];
    assign inter_2[162] = inter_1[162];
    assign inter_2[163] = inter_1[163];
    assign inter_2[164] = inter_1[164]^inter_1[166];
    assign inter_2[165] = inter_1[165]^inter_1[167];
    assign inter_2[166] = inter_1[166];
    assign inter_2[167] = inter_1[167];
    assign inter_2[168] = inter_1[168]^inter_1[170];
    assign inter_2[169] = inter_1[169]^inter_1[171];
    assign inter_2[170] = inter_1[170];
    assign inter_2[171] = inter_1[171];
    assign inter_2[172] = inter_1[172]^inter_1[174];
    assign inter_2[173] = inter_1[173]^inter_1[175];
    assign inter_2[174] = inter_1[174];
    assign inter_2[175] = inter_1[175];
    assign inter_2[176] = inter_1[176]^inter_1[178];
    assign inter_2[177] = inter_1[177]^inter_1[179];
    assign inter_2[178] = inter_1[178];
    assign inter_2[179] = inter_1[179];
    assign inter_2[180] = inter_1[180]^inter_1[182];
    assign inter_2[181] = inter_1[181]^inter_1[183];
    assign inter_2[182] = inter_1[182];
    assign inter_2[183] = inter_1[183];
    assign inter_2[184] = inter_1[184]^inter_1[186];
    assign inter_2[185] = inter_1[185]^inter_1[187];
    assign inter_2[186] = inter_1[186];
    assign inter_2[187] = inter_1[187];
    assign inter_2[188] = inter_1[188]^inter_1[190];
    assign inter_2[189] = inter_1[189]^inter_1[191];
    assign inter_2[190] = inter_1[190];
    assign inter_2[191] = inter_1[191];
    assign inter_2[192] = inter_1[192]^inter_1[194];
    assign inter_2[193] = inter_1[193]^inter_1[195];
    assign inter_2[194] = inter_1[194];
    assign inter_2[195] = inter_1[195];
    assign inter_2[196] = inter_1[196]^inter_1[198];
    assign inter_2[197] = inter_1[197]^inter_1[199];
    assign inter_2[198] = inter_1[198];
    assign inter_2[199] = inter_1[199];
    assign inter_2[200] = inter_1[200]^inter_1[202];
    assign inter_2[201] = inter_1[201]^inter_1[203];
    assign inter_2[202] = inter_1[202];
    assign inter_2[203] = inter_1[203];
    assign inter_2[204] = inter_1[204]^inter_1[206];
    assign inter_2[205] = inter_1[205]^inter_1[207];
    assign inter_2[206] = inter_1[206];
    assign inter_2[207] = inter_1[207];
    assign inter_2[208] = inter_1[208]^inter_1[210];
    assign inter_2[209] = inter_1[209]^inter_1[211];
    assign inter_2[210] = inter_1[210];
    assign inter_2[211] = inter_1[211];
    assign inter_2[212] = inter_1[212]^inter_1[214];
    assign inter_2[213] = inter_1[213]^inter_1[215];
    assign inter_2[214] = inter_1[214];
    assign inter_2[215] = inter_1[215];
    assign inter_2[216] = inter_1[216]^inter_1[218];
    assign inter_2[217] = inter_1[217]^inter_1[219];
    assign inter_2[218] = inter_1[218];
    assign inter_2[219] = inter_1[219];
    assign inter_2[220] = inter_1[220]^inter_1[222];
    assign inter_2[221] = inter_1[221]^inter_1[223];
    assign inter_2[222] = inter_1[222];
    assign inter_2[223] = inter_1[223];
    assign inter_2[224] = inter_1[224]^inter_1[226];
    assign inter_2[225] = inter_1[225]^inter_1[227];
    assign inter_2[226] = inter_1[226];
    assign inter_2[227] = inter_1[227];
    assign inter_2[228] = inter_1[228]^inter_1[230];
    assign inter_2[229] = inter_1[229]^inter_1[231];
    assign inter_2[230] = inter_1[230];
    assign inter_2[231] = inter_1[231];
    assign inter_2[232] = inter_1[232]^inter_1[234];
    assign inter_2[233] = inter_1[233]^inter_1[235];
    assign inter_2[234] = inter_1[234];
    assign inter_2[235] = inter_1[235];
    assign inter_2[236] = inter_1[236]^inter_1[238];
    assign inter_2[237] = inter_1[237]^inter_1[239];
    assign inter_2[238] = inter_1[238];
    assign inter_2[239] = inter_1[239];
    assign inter_2[240] = inter_1[240]^inter_1[242];
    assign inter_2[241] = inter_1[241]^inter_1[243];
    assign inter_2[242] = inter_1[242];
    assign inter_2[243] = inter_1[243];
    assign inter_2[244] = inter_1[244]^inter_1[246];
    assign inter_2[245] = inter_1[245]^inter_1[247];
    assign inter_2[246] = inter_1[246];
    assign inter_2[247] = inter_1[247];
    assign inter_2[248] = inter_1[248]^inter_1[250];
    assign inter_2[249] = inter_1[249]^inter_1[251];
    assign inter_2[250] = inter_1[250];
    assign inter_2[251] = inter_1[251];
    assign inter_2[252] = inter_1[252]^inter_1[254];
    assign inter_2[253] = inter_1[253]^inter_1[255];
    assign inter_2[254] = inter_1[254];
    assign inter_2[255] = inter_1[255];
    assign inter_2[256] = inter_1[256]^inter_1[258];
    assign inter_2[257] = inter_1[257]^inter_1[259];
    assign inter_2[258] = inter_1[258];
    assign inter_2[259] = inter_1[259];
    assign inter_2[260] = inter_1[260]^inter_1[262];
    assign inter_2[261] = inter_1[261]^inter_1[263];
    assign inter_2[262] = inter_1[262];
    assign inter_2[263] = inter_1[263];
    assign inter_2[264] = inter_1[264]^inter_1[266];
    assign inter_2[265] = inter_1[265]^inter_1[267];
    assign inter_2[266] = inter_1[266];
    assign inter_2[267] = inter_1[267];
    assign inter_2[268] = inter_1[268]^inter_1[270];
    assign inter_2[269] = inter_1[269]^inter_1[271];
    assign inter_2[270] = inter_1[270];
    assign inter_2[271] = inter_1[271];
    assign inter_2[272] = inter_1[272]^inter_1[274];
    assign inter_2[273] = inter_1[273]^inter_1[275];
    assign inter_2[274] = inter_1[274];
    assign inter_2[275] = inter_1[275];
    assign inter_2[276] = inter_1[276]^inter_1[278];
    assign inter_2[277] = inter_1[277]^inter_1[279];
    assign inter_2[278] = inter_1[278];
    assign inter_2[279] = inter_1[279];
    assign inter_2[280] = inter_1[280]^inter_1[282];
    assign inter_2[281] = inter_1[281]^inter_1[283];
    assign inter_2[282] = inter_1[282];
    assign inter_2[283] = inter_1[283];
    assign inter_2[284] = inter_1[284]^inter_1[286];
    assign inter_2[285] = inter_1[285]^inter_1[287];
    assign inter_2[286] = inter_1[286];
    assign inter_2[287] = inter_1[287];
    assign inter_2[288] = inter_1[288]^inter_1[290];
    assign inter_2[289] = inter_1[289]^inter_1[291];
    assign inter_2[290] = inter_1[290];
    assign inter_2[291] = inter_1[291];
    assign inter_2[292] = inter_1[292]^inter_1[294];
    assign inter_2[293] = inter_1[293]^inter_1[295];
    assign inter_2[294] = inter_1[294];
    assign inter_2[295] = inter_1[295];
    assign inter_2[296] = inter_1[296]^inter_1[298];
    assign inter_2[297] = inter_1[297]^inter_1[299];
    assign inter_2[298] = inter_1[298];
    assign inter_2[299] = inter_1[299];
    assign inter_2[300] = inter_1[300]^inter_1[302];
    assign inter_2[301] = inter_1[301]^inter_1[303];
    assign inter_2[302] = inter_1[302];
    assign inter_2[303] = inter_1[303];
    assign inter_2[304] = inter_1[304]^inter_1[306];
    assign inter_2[305] = inter_1[305]^inter_1[307];
    assign inter_2[306] = inter_1[306];
    assign inter_2[307] = inter_1[307];
    assign inter_2[308] = inter_1[308]^inter_1[310];
    assign inter_2[309] = inter_1[309]^inter_1[311];
    assign inter_2[310] = inter_1[310];
    assign inter_2[311] = inter_1[311];
    assign inter_2[312] = inter_1[312]^inter_1[314];
    assign inter_2[313] = inter_1[313]^inter_1[315];
    assign inter_2[314] = inter_1[314];
    assign inter_2[315] = inter_1[315];
    assign inter_2[316] = inter_1[316]^inter_1[318];
    assign inter_2[317] = inter_1[317]^inter_1[319];
    assign inter_2[318] = inter_1[318];
    assign inter_2[319] = inter_1[319];
    assign inter_2[320] = inter_1[320]^inter_1[322];
    assign inter_2[321] = inter_1[321]^inter_1[323];
    assign inter_2[322] = inter_1[322];
    assign inter_2[323] = inter_1[323];
    assign inter_2[324] = inter_1[324]^inter_1[326];
    assign inter_2[325] = inter_1[325]^inter_1[327];
    assign inter_2[326] = inter_1[326];
    assign inter_2[327] = inter_1[327];
    assign inter_2[328] = inter_1[328]^inter_1[330];
    assign inter_2[329] = inter_1[329]^inter_1[331];
    assign inter_2[330] = inter_1[330];
    assign inter_2[331] = inter_1[331];
    assign inter_2[332] = inter_1[332]^inter_1[334];
    assign inter_2[333] = inter_1[333]^inter_1[335];
    assign inter_2[334] = inter_1[334];
    assign inter_2[335] = inter_1[335];
    assign inter_2[336] = inter_1[336]^inter_1[338];
    assign inter_2[337] = inter_1[337]^inter_1[339];
    assign inter_2[338] = inter_1[338];
    assign inter_2[339] = inter_1[339];
    assign inter_2[340] = inter_1[340]^inter_1[342];
    assign inter_2[341] = inter_1[341]^inter_1[343];
    assign inter_2[342] = inter_1[342];
    assign inter_2[343] = inter_1[343];
    assign inter_2[344] = inter_1[344]^inter_1[346];
    assign inter_2[345] = inter_1[345]^inter_1[347];
    assign inter_2[346] = inter_1[346];
    assign inter_2[347] = inter_1[347];
    assign inter_2[348] = inter_1[348]^inter_1[350];
    assign inter_2[349] = inter_1[349]^inter_1[351];
    assign inter_2[350] = inter_1[350];
    assign inter_2[351] = inter_1[351];
    assign inter_2[352] = inter_1[352]^inter_1[354];
    assign inter_2[353] = inter_1[353]^inter_1[355];
    assign inter_2[354] = inter_1[354];
    assign inter_2[355] = inter_1[355];
    assign inter_2[356] = inter_1[356]^inter_1[358];
    assign inter_2[357] = inter_1[357]^inter_1[359];
    assign inter_2[358] = inter_1[358];
    assign inter_2[359] = inter_1[359];
    assign inter_2[360] = inter_1[360]^inter_1[362];
    assign inter_2[361] = inter_1[361]^inter_1[363];
    assign inter_2[362] = inter_1[362];
    assign inter_2[363] = inter_1[363];
    assign inter_2[364] = inter_1[364]^inter_1[366];
    assign inter_2[365] = inter_1[365]^inter_1[367];
    assign inter_2[366] = inter_1[366];
    assign inter_2[367] = inter_1[367];
    assign inter_2[368] = inter_1[368]^inter_1[370];
    assign inter_2[369] = inter_1[369]^inter_1[371];
    assign inter_2[370] = inter_1[370];
    assign inter_2[371] = inter_1[371];
    assign inter_2[372] = inter_1[372]^inter_1[374];
    assign inter_2[373] = inter_1[373]^inter_1[375];
    assign inter_2[374] = inter_1[374];
    assign inter_2[375] = inter_1[375];
    assign inter_2[376] = inter_1[376]^inter_1[378];
    assign inter_2[377] = inter_1[377]^inter_1[379];
    assign inter_2[378] = inter_1[378];
    assign inter_2[379] = inter_1[379];
    assign inter_2[380] = inter_1[380]^inter_1[382];
    assign inter_2[381] = inter_1[381]^inter_1[383];
    assign inter_2[382] = inter_1[382];
    assign inter_2[383] = inter_1[383];
    assign inter_2[384] = inter_1[384]^inter_1[386];
    assign inter_2[385] = inter_1[385]^inter_1[387];
    assign inter_2[386] = inter_1[386];
    assign inter_2[387] = inter_1[387];
    assign inter_2[388] = inter_1[388]^inter_1[390];
    assign inter_2[389] = inter_1[389]^inter_1[391];
    assign inter_2[390] = inter_1[390];
    assign inter_2[391] = inter_1[391];
    assign inter_2[392] = inter_1[392]^inter_1[394];
    assign inter_2[393] = inter_1[393]^inter_1[395];
    assign inter_2[394] = inter_1[394];
    assign inter_2[395] = inter_1[395];
    assign inter_2[396] = inter_1[396]^inter_1[398];
    assign inter_2[397] = inter_1[397]^inter_1[399];
    assign inter_2[398] = inter_1[398];
    assign inter_2[399] = inter_1[399];
    assign inter_2[400] = inter_1[400]^inter_1[402];
    assign inter_2[401] = inter_1[401]^inter_1[403];
    assign inter_2[402] = inter_1[402];
    assign inter_2[403] = inter_1[403];
    assign inter_2[404] = inter_1[404]^inter_1[406];
    assign inter_2[405] = inter_1[405]^inter_1[407];
    assign inter_2[406] = inter_1[406];
    assign inter_2[407] = inter_1[407];
    assign inter_2[408] = inter_1[408]^inter_1[410];
    assign inter_2[409] = inter_1[409]^inter_1[411];
    assign inter_2[410] = inter_1[410];
    assign inter_2[411] = inter_1[411];
    assign inter_2[412] = inter_1[412]^inter_1[414];
    assign inter_2[413] = inter_1[413]^inter_1[415];
    assign inter_2[414] = inter_1[414];
    assign inter_2[415] = inter_1[415];
    assign inter_2[416] = inter_1[416]^inter_1[418];
    assign inter_2[417] = inter_1[417]^inter_1[419];
    assign inter_2[418] = inter_1[418];
    assign inter_2[419] = inter_1[419];
    assign inter_2[420] = inter_1[420]^inter_1[422];
    assign inter_2[421] = inter_1[421]^inter_1[423];
    assign inter_2[422] = inter_1[422];
    assign inter_2[423] = inter_1[423];
    assign inter_2[424] = inter_1[424]^inter_1[426];
    assign inter_2[425] = inter_1[425]^inter_1[427];
    assign inter_2[426] = inter_1[426];
    assign inter_2[427] = inter_1[427];
    assign inter_2[428] = inter_1[428]^inter_1[430];
    assign inter_2[429] = inter_1[429]^inter_1[431];
    assign inter_2[430] = inter_1[430];
    assign inter_2[431] = inter_1[431];
    assign inter_2[432] = inter_1[432]^inter_1[434];
    assign inter_2[433] = inter_1[433]^inter_1[435];
    assign inter_2[434] = inter_1[434];
    assign inter_2[435] = inter_1[435];
    assign inter_2[436] = inter_1[436]^inter_1[438];
    assign inter_2[437] = inter_1[437]^inter_1[439];
    assign inter_2[438] = inter_1[438];
    assign inter_2[439] = inter_1[439];
    assign inter_2[440] = inter_1[440]^inter_1[442];
    assign inter_2[441] = inter_1[441]^inter_1[443];
    assign inter_2[442] = inter_1[442];
    assign inter_2[443] = inter_1[443];
    assign inter_2[444] = inter_1[444]^inter_1[446];
    assign inter_2[445] = inter_1[445]^inter_1[447];
    assign inter_2[446] = inter_1[446];
    assign inter_2[447] = inter_1[447];
    assign inter_2[448] = inter_1[448]^inter_1[450];
    assign inter_2[449] = inter_1[449]^inter_1[451];
    assign inter_2[450] = inter_1[450];
    assign inter_2[451] = inter_1[451];
    assign inter_2[452] = inter_1[452]^inter_1[454];
    assign inter_2[453] = inter_1[453]^inter_1[455];
    assign inter_2[454] = inter_1[454];
    assign inter_2[455] = inter_1[455];
    assign inter_2[456] = inter_1[456]^inter_1[458];
    assign inter_2[457] = inter_1[457]^inter_1[459];
    assign inter_2[458] = inter_1[458];
    assign inter_2[459] = inter_1[459];
    assign inter_2[460] = inter_1[460]^inter_1[462];
    assign inter_2[461] = inter_1[461]^inter_1[463];
    assign inter_2[462] = inter_1[462];
    assign inter_2[463] = inter_1[463];
    assign inter_2[464] = inter_1[464]^inter_1[466];
    assign inter_2[465] = inter_1[465]^inter_1[467];
    assign inter_2[466] = inter_1[466];
    assign inter_2[467] = inter_1[467];
    assign inter_2[468] = inter_1[468]^inter_1[470];
    assign inter_2[469] = inter_1[469]^inter_1[471];
    assign inter_2[470] = inter_1[470];
    assign inter_2[471] = inter_1[471];
    assign inter_2[472] = inter_1[472]^inter_1[474];
    assign inter_2[473] = inter_1[473]^inter_1[475];
    assign inter_2[474] = inter_1[474];
    assign inter_2[475] = inter_1[475];
    assign inter_2[476] = inter_1[476]^inter_1[478];
    assign inter_2[477] = inter_1[477]^inter_1[479];
    assign inter_2[478] = inter_1[478];
    assign inter_2[479] = inter_1[479];
    assign inter_2[480] = inter_1[480]^inter_1[482];
    assign inter_2[481] = inter_1[481]^inter_1[483];
    assign inter_2[482] = inter_1[482];
    assign inter_2[483] = inter_1[483];
    assign inter_2[484] = inter_1[484]^inter_1[486];
    assign inter_2[485] = inter_1[485]^inter_1[487];
    assign inter_2[486] = inter_1[486];
    assign inter_2[487] = inter_1[487];
    assign inter_2[488] = inter_1[488]^inter_1[490];
    assign inter_2[489] = inter_1[489]^inter_1[491];
    assign inter_2[490] = inter_1[490];
    assign inter_2[491] = inter_1[491];
    assign inter_2[492] = inter_1[492]^inter_1[494];
    assign inter_2[493] = inter_1[493]^inter_1[495];
    assign inter_2[494] = inter_1[494];
    assign inter_2[495] = inter_1[495];
    assign inter_2[496] = inter_1[496]^inter_1[498];
    assign inter_2[497] = inter_1[497]^inter_1[499];
    assign inter_2[498] = inter_1[498];
    assign inter_2[499] = inter_1[499];
    assign inter_2[500] = inter_1[500]^inter_1[502];
    assign inter_2[501] = inter_1[501]^inter_1[503];
    assign inter_2[502] = inter_1[502];
    assign inter_2[503] = inter_1[503];
    assign inter_2[504] = inter_1[504]^inter_1[506];
    assign inter_2[505] = inter_1[505]^inter_1[507];
    assign inter_2[506] = inter_1[506];
    assign inter_2[507] = inter_1[507];
    assign inter_2[508] = inter_1[508]^inter_1[510];
    assign inter_2[509] = inter_1[509]^inter_1[511];
    assign inter_2[510] = inter_1[510];
    assign inter_2[511] = inter_1[511];
    assign inter_2[512] = inter_1[512]^inter_1[514];
    assign inter_2[513] = inter_1[513]^inter_1[515];
    assign inter_2[514] = inter_1[514];
    assign inter_2[515] = inter_1[515];
    assign inter_2[516] = inter_1[516]^inter_1[518];
    assign inter_2[517] = inter_1[517]^inter_1[519];
    assign inter_2[518] = inter_1[518];
    assign inter_2[519] = inter_1[519];
    assign inter_2[520] = inter_1[520]^inter_1[522];
    assign inter_2[521] = inter_1[521]^inter_1[523];
    assign inter_2[522] = inter_1[522];
    assign inter_2[523] = inter_1[523];
    assign inter_2[524] = inter_1[524]^inter_1[526];
    assign inter_2[525] = inter_1[525]^inter_1[527];
    assign inter_2[526] = inter_1[526];
    assign inter_2[527] = inter_1[527];
    assign inter_2[528] = inter_1[528]^inter_1[530];
    assign inter_2[529] = inter_1[529]^inter_1[531];
    assign inter_2[530] = inter_1[530];
    assign inter_2[531] = inter_1[531];
    assign inter_2[532] = inter_1[532]^inter_1[534];
    assign inter_2[533] = inter_1[533]^inter_1[535];
    assign inter_2[534] = inter_1[534];
    assign inter_2[535] = inter_1[535];
    assign inter_2[536] = inter_1[536]^inter_1[538];
    assign inter_2[537] = inter_1[537]^inter_1[539];
    assign inter_2[538] = inter_1[538];
    assign inter_2[539] = inter_1[539];
    assign inter_2[540] = inter_1[540]^inter_1[542];
    assign inter_2[541] = inter_1[541]^inter_1[543];
    assign inter_2[542] = inter_1[542];
    assign inter_2[543] = inter_1[543];
    assign inter_2[544] = inter_1[544]^inter_1[546];
    assign inter_2[545] = inter_1[545]^inter_1[547];
    assign inter_2[546] = inter_1[546];
    assign inter_2[547] = inter_1[547];
    assign inter_2[548] = inter_1[548]^inter_1[550];
    assign inter_2[549] = inter_1[549]^inter_1[551];
    assign inter_2[550] = inter_1[550];
    assign inter_2[551] = inter_1[551];
    assign inter_2[552] = inter_1[552]^inter_1[554];
    assign inter_2[553] = inter_1[553]^inter_1[555];
    assign inter_2[554] = inter_1[554];
    assign inter_2[555] = inter_1[555];
    assign inter_2[556] = inter_1[556]^inter_1[558];
    assign inter_2[557] = inter_1[557]^inter_1[559];
    assign inter_2[558] = inter_1[558];
    assign inter_2[559] = inter_1[559];
    assign inter_2[560] = inter_1[560]^inter_1[562];
    assign inter_2[561] = inter_1[561]^inter_1[563];
    assign inter_2[562] = inter_1[562];
    assign inter_2[563] = inter_1[563];
    assign inter_2[564] = inter_1[564]^inter_1[566];
    assign inter_2[565] = inter_1[565]^inter_1[567];
    assign inter_2[566] = inter_1[566];
    assign inter_2[567] = inter_1[567];
    assign inter_2[568] = inter_1[568]^inter_1[570];
    assign inter_2[569] = inter_1[569]^inter_1[571];
    assign inter_2[570] = inter_1[570];
    assign inter_2[571] = inter_1[571];
    assign inter_2[572] = inter_1[572]^inter_1[574];
    assign inter_2[573] = inter_1[573]^inter_1[575];
    assign inter_2[574] = inter_1[574];
    assign inter_2[575] = inter_1[575];
    assign inter_2[576] = inter_1[576]^inter_1[578];
    assign inter_2[577] = inter_1[577]^inter_1[579];
    assign inter_2[578] = inter_1[578];
    assign inter_2[579] = inter_1[579];
    assign inter_2[580] = inter_1[580]^inter_1[582];
    assign inter_2[581] = inter_1[581]^inter_1[583];
    assign inter_2[582] = inter_1[582];
    assign inter_2[583] = inter_1[583];
    assign inter_2[584] = inter_1[584]^inter_1[586];
    assign inter_2[585] = inter_1[585]^inter_1[587];
    assign inter_2[586] = inter_1[586];
    assign inter_2[587] = inter_1[587];
    assign inter_2[588] = inter_1[588]^inter_1[590];
    assign inter_2[589] = inter_1[589]^inter_1[591];
    assign inter_2[590] = inter_1[590];
    assign inter_2[591] = inter_1[591];
    assign inter_2[592] = inter_1[592]^inter_1[594];
    assign inter_2[593] = inter_1[593]^inter_1[595];
    assign inter_2[594] = inter_1[594];
    assign inter_2[595] = inter_1[595];
    assign inter_2[596] = inter_1[596]^inter_1[598];
    assign inter_2[597] = inter_1[597]^inter_1[599];
    assign inter_2[598] = inter_1[598];
    assign inter_2[599] = inter_1[599];
    assign inter_2[600] = inter_1[600]^inter_1[602];
    assign inter_2[601] = inter_1[601]^inter_1[603];
    assign inter_2[602] = inter_1[602];
    assign inter_2[603] = inter_1[603];
    assign inter_2[604] = inter_1[604]^inter_1[606];
    assign inter_2[605] = inter_1[605]^inter_1[607];
    assign inter_2[606] = inter_1[606];
    assign inter_2[607] = inter_1[607];
    assign inter_2[608] = inter_1[608]^inter_1[610];
    assign inter_2[609] = inter_1[609]^inter_1[611];
    assign inter_2[610] = inter_1[610];
    assign inter_2[611] = inter_1[611];
    assign inter_2[612] = inter_1[612]^inter_1[614];
    assign inter_2[613] = inter_1[613]^inter_1[615];
    assign inter_2[614] = inter_1[614];
    assign inter_2[615] = inter_1[615];
    assign inter_2[616] = inter_1[616]^inter_1[618];
    assign inter_2[617] = inter_1[617]^inter_1[619];
    assign inter_2[618] = inter_1[618];
    assign inter_2[619] = inter_1[619];
    assign inter_2[620] = inter_1[620]^inter_1[622];
    assign inter_2[621] = inter_1[621]^inter_1[623];
    assign inter_2[622] = inter_1[622];
    assign inter_2[623] = inter_1[623];
    assign inter_2[624] = inter_1[624]^inter_1[626];
    assign inter_2[625] = inter_1[625]^inter_1[627];
    assign inter_2[626] = inter_1[626];
    assign inter_2[627] = inter_1[627];
    assign inter_2[628] = inter_1[628]^inter_1[630];
    assign inter_2[629] = inter_1[629]^inter_1[631];
    assign inter_2[630] = inter_1[630];
    assign inter_2[631] = inter_1[631];
    assign inter_2[632] = inter_1[632]^inter_1[634];
    assign inter_2[633] = inter_1[633]^inter_1[635];
    assign inter_2[634] = inter_1[634];
    assign inter_2[635] = inter_1[635];
    assign inter_2[636] = inter_1[636]^inter_1[638];
    assign inter_2[637] = inter_1[637]^inter_1[639];
    assign inter_2[638] = inter_1[638];
    assign inter_2[639] = inter_1[639];
    assign inter_2[640] = inter_1[640]^inter_1[642];
    assign inter_2[641] = inter_1[641]^inter_1[643];
    assign inter_2[642] = inter_1[642];
    assign inter_2[643] = inter_1[643];
    assign inter_2[644] = inter_1[644]^inter_1[646];
    assign inter_2[645] = inter_1[645]^inter_1[647];
    assign inter_2[646] = inter_1[646];
    assign inter_2[647] = inter_1[647];
    assign inter_2[648] = inter_1[648]^inter_1[650];
    assign inter_2[649] = inter_1[649]^inter_1[651];
    assign inter_2[650] = inter_1[650];
    assign inter_2[651] = inter_1[651];
    assign inter_2[652] = inter_1[652]^inter_1[654];
    assign inter_2[653] = inter_1[653]^inter_1[655];
    assign inter_2[654] = inter_1[654];
    assign inter_2[655] = inter_1[655];
    assign inter_2[656] = inter_1[656]^inter_1[658];
    assign inter_2[657] = inter_1[657]^inter_1[659];
    assign inter_2[658] = inter_1[658];
    assign inter_2[659] = inter_1[659];
    assign inter_2[660] = inter_1[660]^inter_1[662];
    assign inter_2[661] = inter_1[661]^inter_1[663];
    assign inter_2[662] = inter_1[662];
    assign inter_2[663] = inter_1[663];
    assign inter_2[664] = inter_1[664]^inter_1[666];
    assign inter_2[665] = inter_1[665]^inter_1[667];
    assign inter_2[666] = inter_1[666];
    assign inter_2[667] = inter_1[667];
    assign inter_2[668] = inter_1[668]^inter_1[670];
    assign inter_2[669] = inter_1[669]^inter_1[671];
    assign inter_2[670] = inter_1[670];
    assign inter_2[671] = inter_1[671];
    assign inter_2[672] = inter_1[672]^inter_1[674];
    assign inter_2[673] = inter_1[673]^inter_1[675];
    assign inter_2[674] = inter_1[674];
    assign inter_2[675] = inter_1[675];
    assign inter_2[676] = inter_1[676]^inter_1[678];
    assign inter_2[677] = inter_1[677]^inter_1[679];
    assign inter_2[678] = inter_1[678];
    assign inter_2[679] = inter_1[679];
    assign inter_2[680] = inter_1[680]^inter_1[682];
    assign inter_2[681] = inter_1[681]^inter_1[683];
    assign inter_2[682] = inter_1[682];
    assign inter_2[683] = inter_1[683];
    assign inter_2[684] = inter_1[684]^inter_1[686];
    assign inter_2[685] = inter_1[685]^inter_1[687];
    assign inter_2[686] = inter_1[686];
    assign inter_2[687] = inter_1[687];
    assign inter_2[688] = inter_1[688]^inter_1[690];
    assign inter_2[689] = inter_1[689]^inter_1[691];
    assign inter_2[690] = inter_1[690];
    assign inter_2[691] = inter_1[691];
    assign inter_2[692] = inter_1[692]^inter_1[694];
    assign inter_2[693] = inter_1[693]^inter_1[695];
    assign inter_2[694] = inter_1[694];
    assign inter_2[695] = inter_1[695];
    assign inter_2[696] = inter_1[696]^inter_1[698];
    assign inter_2[697] = inter_1[697]^inter_1[699];
    assign inter_2[698] = inter_1[698];
    assign inter_2[699] = inter_1[699];
    assign inter_2[700] = inter_1[700]^inter_1[702];
    assign inter_2[701] = inter_1[701]^inter_1[703];
    assign inter_2[702] = inter_1[702];
    assign inter_2[703] = inter_1[703];
    assign inter_2[704] = inter_1[704]^inter_1[706];
    assign inter_2[705] = inter_1[705]^inter_1[707];
    assign inter_2[706] = inter_1[706];
    assign inter_2[707] = inter_1[707];
    assign inter_2[708] = inter_1[708]^inter_1[710];
    assign inter_2[709] = inter_1[709]^inter_1[711];
    assign inter_2[710] = inter_1[710];
    assign inter_2[711] = inter_1[711];
    assign inter_2[712] = inter_1[712]^inter_1[714];
    assign inter_2[713] = inter_1[713]^inter_1[715];
    assign inter_2[714] = inter_1[714];
    assign inter_2[715] = inter_1[715];
    assign inter_2[716] = inter_1[716]^inter_1[718];
    assign inter_2[717] = inter_1[717]^inter_1[719];
    assign inter_2[718] = inter_1[718];
    assign inter_2[719] = inter_1[719];
    assign inter_2[720] = inter_1[720]^inter_1[722];
    assign inter_2[721] = inter_1[721]^inter_1[723];
    assign inter_2[722] = inter_1[722];
    assign inter_2[723] = inter_1[723];
    assign inter_2[724] = inter_1[724]^inter_1[726];
    assign inter_2[725] = inter_1[725]^inter_1[727];
    assign inter_2[726] = inter_1[726];
    assign inter_2[727] = inter_1[727];
    assign inter_2[728] = inter_1[728]^inter_1[730];
    assign inter_2[729] = inter_1[729]^inter_1[731];
    assign inter_2[730] = inter_1[730];
    assign inter_2[731] = inter_1[731];
    assign inter_2[732] = inter_1[732]^inter_1[734];
    assign inter_2[733] = inter_1[733]^inter_1[735];
    assign inter_2[734] = inter_1[734];
    assign inter_2[735] = inter_1[735];
    assign inter_2[736] = inter_1[736]^inter_1[738];
    assign inter_2[737] = inter_1[737]^inter_1[739];
    assign inter_2[738] = inter_1[738];
    assign inter_2[739] = inter_1[739];
    assign inter_2[740] = inter_1[740]^inter_1[742];
    assign inter_2[741] = inter_1[741]^inter_1[743];
    assign inter_2[742] = inter_1[742];
    assign inter_2[743] = inter_1[743];
    assign inter_2[744] = inter_1[744]^inter_1[746];
    assign inter_2[745] = inter_1[745]^inter_1[747];
    assign inter_2[746] = inter_1[746];
    assign inter_2[747] = inter_1[747];
    assign inter_2[748] = inter_1[748]^inter_1[750];
    assign inter_2[749] = inter_1[749]^inter_1[751];
    assign inter_2[750] = inter_1[750];
    assign inter_2[751] = inter_1[751];
    assign inter_2[752] = inter_1[752]^inter_1[754];
    assign inter_2[753] = inter_1[753]^inter_1[755];
    assign inter_2[754] = inter_1[754];
    assign inter_2[755] = inter_1[755];
    assign inter_2[756] = inter_1[756]^inter_1[758];
    assign inter_2[757] = inter_1[757]^inter_1[759];
    assign inter_2[758] = inter_1[758];
    assign inter_2[759] = inter_1[759];
    assign inter_2[760] = inter_1[760]^inter_1[762];
    assign inter_2[761] = inter_1[761]^inter_1[763];
    assign inter_2[762] = inter_1[762];
    assign inter_2[763] = inter_1[763];
    assign inter_2[764] = inter_1[764]^inter_1[766];
    assign inter_2[765] = inter_1[765]^inter_1[767];
    assign inter_2[766] = inter_1[766];
    assign inter_2[767] = inter_1[767];
    assign inter_2[768] = inter_1[768]^inter_1[770];
    assign inter_2[769] = inter_1[769]^inter_1[771];
    assign inter_2[770] = inter_1[770];
    assign inter_2[771] = inter_1[771];
    assign inter_2[772] = inter_1[772]^inter_1[774];
    assign inter_2[773] = inter_1[773]^inter_1[775];
    assign inter_2[774] = inter_1[774];
    assign inter_2[775] = inter_1[775];
    assign inter_2[776] = inter_1[776]^inter_1[778];
    assign inter_2[777] = inter_1[777]^inter_1[779];
    assign inter_2[778] = inter_1[778];
    assign inter_2[779] = inter_1[779];
    assign inter_2[780] = inter_1[780]^inter_1[782];
    assign inter_2[781] = inter_1[781]^inter_1[783];
    assign inter_2[782] = inter_1[782];
    assign inter_2[783] = inter_1[783];
    assign inter_2[784] = inter_1[784]^inter_1[786];
    assign inter_2[785] = inter_1[785]^inter_1[787];
    assign inter_2[786] = inter_1[786];
    assign inter_2[787] = inter_1[787];
    assign inter_2[788] = inter_1[788]^inter_1[790];
    assign inter_2[789] = inter_1[789]^inter_1[791];
    assign inter_2[790] = inter_1[790];
    assign inter_2[791] = inter_1[791];
    assign inter_2[792] = inter_1[792]^inter_1[794];
    assign inter_2[793] = inter_1[793]^inter_1[795];
    assign inter_2[794] = inter_1[794];
    assign inter_2[795] = inter_1[795];
    assign inter_2[796] = inter_1[796]^inter_1[798];
    assign inter_2[797] = inter_1[797]^inter_1[799];
    assign inter_2[798] = inter_1[798];
    assign inter_2[799] = inter_1[799];
    assign inter_2[800] = inter_1[800]^inter_1[802];
    assign inter_2[801] = inter_1[801]^inter_1[803];
    assign inter_2[802] = inter_1[802];
    assign inter_2[803] = inter_1[803];
    assign inter_2[804] = inter_1[804]^inter_1[806];
    assign inter_2[805] = inter_1[805]^inter_1[807];
    assign inter_2[806] = inter_1[806];
    assign inter_2[807] = inter_1[807];
    assign inter_2[808] = inter_1[808]^inter_1[810];
    assign inter_2[809] = inter_1[809]^inter_1[811];
    assign inter_2[810] = inter_1[810];
    assign inter_2[811] = inter_1[811];
    assign inter_2[812] = inter_1[812]^inter_1[814];
    assign inter_2[813] = inter_1[813]^inter_1[815];
    assign inter_2[814] = inter_1[814];
    assign inter_2[815] = inter_1[815];
    assign inter_2[816] = inter_1[816]^inter_1[818];
    assign inter_2[817] = inter_1[817]^inter_1[819];
    assign inter_2[818] = inter_1[818];
    assign inter_2[819] = inter_1[819];
    assign inter_2[820] = inter_1[820]^inter_1[822];
    assign inter_2[821] = inter_1[821]^inter_1[823];
    assign inter_2[822] = inter_1[822];
    assign inter_2[823] = inter_1[823];
    assign inter_2[824] = inter_1[824]^inter_1[826];
    assign inter_2[825] = inter_1[825]^inter_1[827];
    assign inter_2[826] = inter_1[826];
    assign inter_2[827] = inter_1[827];
    assign inter_2[828] = inter_1[828]^inter_1[830];
    assign inter_2[829] = inter_1[829]^inter_1[831];
    assign inter_2[830] = inter_1[830];
    assign inter_2[831] = inter_1[831];
    assign inter_2[832] = inter_1[832]^inter_1[834];
    assign inter_2[833] = inter_1[833]^inter_1[835];
    assign inter_2[834] = inter_1[834];
    assign inter_2[835] = inter_1[835];
    assign inter_2[836] = inter_1[836]^inter_1[838];
    assign inter_2[837] = inter_1[837]^inter_1[839];
    assign inter_2[838] = inter_1[838];
    assign inter_2[839] = inter_1[839];
    assign inter_2[840] = inter_1[840]^inter_1[842];
    assign inter_2[841] = inter_1[841]^inter_1[843];
    assign inter_2[842] = inter_1[842];
    assign inter_2[843] = inter_1[843];
    assign inter_2[844] = inter_1[844]^inter_1[846];
    assign inter_2[845] = inter_1[845]^inter_1[847];
    assign inter_2[846] = inter_1[846];
    assign inter_2[847] = inter_1[847];
    assign inter_2[848] = inter_1[848]^inter_1[850];
    assign inter_2[849] = inter_1[849]^inter_1[851];
    assign inter_2[850] = inter_1[850];
    assign inter_2[851] = inter_1[851];
    assign inter_2[852] = inter_1[852]^inter_1[854];
    assign inter_2[853] = inter_1[853]^inter_1[855];
    assign inter_2[854] = inter_1[854];
    assign inter_2[855] = inter_1[855];
    assign inter_2[856] = inter_1[856]^inter_1[858];
    assign inter_2[857] = inter_1[857]^inter_1[859];
    assign inter_2[858] = inter_1[858];
    assign inter_2[859] = inter_1[859];
    assign inter_2[860] = inter_1[860]^inter_1[862];
    assign inter_2[861] = inter_1[861]^inter_1[863];
    assign inter_2[862] = inter_1[862];
    assign inter_2[863] = inter_1[863];
    assign inter_2[864] = inter_1[864]^inter_1[866];
    assign inter_2[865] = inter_1[865]^inter_1[867];
    assign inter_2[866] = inter_1[866];
    assign inter_2[867] = inter_1[867];
    assign inter_2[868] = inter_1[868]^inter_1[870];
    assign inter_2[869] = inter_1[869]^inter_1[871];
    assign inter_2[870] = inter_1[870];
    assign inter_2[871] = inter_1[871];
    assign inter_2[872] = inter_1[872]^inter_1[874];
    assign inter_2[873] = inter_1[873]^inter_1[875];
    assign inter_2[874] = inter_1[874];
    assign inter_2[875] = inter_1[875];
    assign inter_2[876] = inter_1[876]^inter_1[878];
    assign inter_2[877] = inter_1[877]^inter_1[879];
    assign inter_2[878] = inter_1[878];
    assign inter_2[879] = inter_1[879];
    assign inter_2[880] = inter_1[880]^inter_1[882];
    assign inter_2[881] = inter_1[881]^inter_1[883];
    assign inter_2[882] = inter_1[882];
    assign inter_2[883] = inter_1[883];
    assign inter_2[884] = inter_1[884]^inter_1[886];
    assign inter_2[885] = inter_1[885]^inter_1[887];
    assign inter_2[886] = inter_1[886];
    assign inter_2[887] = inter_1[887];
    assign inter_2[888] = inter_1[888]^inter_1[890];
    assign inter_2[889] = inter_1[889]^inter_1[891];
    assign inter_2[890] = inter_1[890];
    assign inter_2[891] = inter_1[891];
    assign inter_2[892] = inter_1[892]^inter_1[894];
    assign inter_2[893] = inter_1[893]^inter_1[895];
    assign inter_2[894] = inter_1[894];
    assign inter_2[895] = inter_1[895];
    assign inter_2[896] = inter_1[896]^inter_1[898];
    assign inter_2[897] = inter_1[897]^inter_1[899];
    assign inter_2[898] = inter_1[898];
    assign inter_2[899] = inter_1[899];
    assign inter_2[900] = inter_1[900]^inter_1[902];
    assign inter_2[901] = inter_1[901]^inter_1[903];
    assign inter_2[902] = inter_1[902];
    assign inter_2[903] = inter_1[903];
    assign inter_2[904] = inter_1[904]^inter_1[906];
    assign inter_2[905] = inter_1[905]^inter_1[907];
    assign inter_2[906] = inter_1[906];
    assign inter_2[907] = inter_1[907];
    assign inter_2[908] = inter_1[908]^inter_1[910];
    assign inter_2[909] = inter_1[909]^inter_1[911];
    assign inter_2[910] = inter_1[910];
    assign inter_2[911] = inter_1[911];
    assign inter_2[912] = inter_1[912]^inter_1[914];
    assign inter_2[913] = inter_1[913]^inter_1[915];
    assign inter_2[914] = inter_1[914];
    assign inter_2[915] = inter_1[915];
    assign inter_2[916] = inter_1[916]^inter_1[918];
    assign inter_2[917] = inter_1[917]^inter_1[919];
    assign inter_2[918] = inter_1[918];
    assign inter_2[919] = inter_1[919];
    assign inter_2[920] = inter_1[920]^inter_1[922];
    assign inter_2[921] = inter_1[921]^inter_1[923];
    assign inter_2[922] = inter_1[922];
    assign inter_2[923] = inter_1[923];
    assign inter_2[924] = inter_1[924]^inter_1[926];
    assign inter_2[925] = inter_1[925]^inter_1[927];
    assign inter_2[926] = inter_1[926];
    assign inter_2[927] = inter_1[927];
    assign inter_2[928] = inter_1[928]^inter_1[930];
    assign inter_2[929] = inter_1[929]^inter_1[931];
    assign inter_2[930] = inter_1[930];
    assign inter_2[931] = inter_1[931];
    assign inter_2[932] = inter_1[932]^inter_1[934];
    assign inter_2[933] = inter_1[933]^inter_1[935];
    assign inter_2[934] = inter_1[934];
    assign inter_2[935] = inter_1[935];
    assign inter_2[936] = inter_1[936]^inter_1[938];
    assign inter_2[937] = inter_1[937]^inter_1[939];
    assign inter_2[938] = inter_1[938];
    assign inter_2[939] = inter_1[939];
    assign inter_2[940] = inter_1[940]^inter_1[942];
    assign inter_2[941] = inter_1[941]^inter_1[943];
    assign inter_2[942] = inter_1[942];
    assign inter_2[943] = inter_1[943];
    assign inter_2[944] = inter_1[944]^inter_1[946];
    assign inter_2[945] = inter_1[945]^inter_1[947];
    assign inter_2[946] = inter_1[946];
    assign inter_2[947] = inter_1[947];
    assign inter_2[948] = inter_1[948]^inter_1[950];
    assign inter_2[949] = inter_1[949]^inter_1[951];
    assign inter_2[950] = inter_1[950];
    assign inter_2[951] = inter_1[951];
    assign inter_2[952] = inter_1[952]^inter_1[954];
    assign inter_2[953] = inter_1[953]^inter_1[955];
    assign inter_2[954] = inter_1[954];
    assign inter_2[955] = inter_1[955];
    assign inter_2[956] = inter_1[956]^inter_1[958];
    assign inter_2[957] = inter_1[957]^inter_1[959];
    assign inter_2[958] = inter_1[958];
    assign inter_2[959] = inter_1[959];
    assign inter_2[960] = inter_1[960]^inter_1[962];
    assign inter_2[961] = inter_1[961]^inter_1[963];
    assign inter_2[962] = inter_1[962];
    assign inter_2[963] = inter_1[963];
    assign inter_2[964] = inter_1[964]^inter_1[966];
    assign inter_2[965] = inter_1[965]^inter_1[967];
    assign inter_2[966] = inter_1[966];
    assign inter_2[967] = inter_1[967];
    assign inter_2[968] = inter_1[968]^inter_1[970];
    assign inter_2[969] = inter_1[969]^inter_1[971];
    assign inter_2[970] = inter_1[970];
    assign inter_2[971] = inter_1[971];
    assign inter_2[972] = inter_1[972]^inter_1[974];
    assign inter_2[973] = inter_1[973]^inter_1[975];
    assign inter_2[974] = inter_1[974];
    assign inter_2[975] = inter_1[975];
    assign inter_2[976] = inter_1[976]^inter_1[978];
    assign inter_2[977] = inter_1[977]^inter_1[979];
    assign inter_2[978] = inter_1[978];
    assign inter_2[979] = inter_1[979];
    assign inter_2[980] = inter_1[980]^inter_1[982];
    assign inter_2[981] = inter_1[981]^inter_1[983];
    assign inter_2[982] = inter_1[982];
    assign inter_2[983] = inter_1[983];
    assign inter_2[984] = inter_1[984]^inter_1[986];
    assign inter_2[985] = inter_1[985]^inter_1[987];
    assign inter_2[986] = inter_1[986];
    assign inter_2[987] = inter_1[987];
    assign inter_2[988] = inter_1[988]^inter_1[990];
    assign inter_2[989] = inter_1[989]^inter_1[991];
    assign inter_2[990] = inter_1[990];
    assign inter_2[991] = inter_1[991];
    assign inter_2[992] = inter_1[992]^inter_1[994];
    assign inter_2[993] = inter_1[993]^inter_1[995];
    assign inter_2[994] = inter_1[994];
    assign inter_2[995] = inter_1[995];
    assign inter_2[996] = inter_1[996]^inter_1[998];
    assign inter_2[997] = inter_1[997]^inter_1[999];
    assign inter_2[998] = inter_1[998];
    assign inter_2[999] = inter_1[999];
    assign inter_2[1000] = inter_1[1000]^inter_1[1002];
    assign inter_2[1001] = inter_1[1001]^inter_1[1003];
    assign inter_2[1002] = inter_1[1002];
    assign inter_2[1003] = inter_1[1003];
    assign inter_2[1004] = inter_1[1004]^inter_1[1006];
    assign inter_2[1005] = inter_1[1005]^inter_1[1007];
    assign inter_2[1006] = inter_1[1006];
    assign inter_2[1007] = inter_1[1007];
    assign inter_2[1008] = inter_1[1008]^inter_1[1010];
    assign inter_2[1009] = inter_1[1009]^inter_1[1011];
    assign inter_2[1010] = inter_1[1010];
    assign inter_2[1011] = inter_1[1011];
    assign inter_2[1012] = inter_1[1012]^inter_1[1014];
    assign inter_2[1013] = inter_1[1013]^inter_1[1015];
    assign inter_2[1014] = inter_1[1014];
    assign inter_2[1015] = inter_1[1015];
    assign inter_2[1016] = inter_1[1016]^inter_1[1018];
    assign inter_2[1017] = inter_1[1017]^inter_1[1019];
    assign inter_2[1018] = inter_1[1018];
    assign inter_2[1019] = inter_1[1019];
    assign inter_2[1020] = inter_1[1020]^inter_1[1022];
    assign inter_2[1021] = inter_1[1021]^inter_1[1023];
    assign inter_2[1022] = inter_1[1022];
    assign inter_2[1023] = inter_1[1023];
    /***************************/
    assign inter_3[0] = inter_2[0]^inter_2[4];
    assign inter_3[1] = inter_2[1]^inter_2[5];
    assign inter_3[2] = inter_2[2]^inter_2[6];
    assign inter_3[3] = inter_2[3]^inter_2[7];
    assign inter_3[4] = inter_2[4];
    assign inter_3[5] = inter_2[5];
    assign inter_3[6] = inter_2[6];
    assign inter_3[7] = inter_2[7];
    assign inter_3[8] = inter_2[8]^inter_2[12];
    assign inter_3[9] = inter_2[9]^inter_2[13];
    assign inter_3[10] = inter_2[10]^inter_2[14];
    assign inter_3[11] = inter_2[11]^inter_2[15];
    assign inter_3[12] = inter_2[12];
    assign inter_3[13] = inter_2[13];
    assign inter_3[14] = inter_2[14];
    assign inter_3[15] = inter_2[15];
    assign inter_3[16] = inter_2[16]^inter_2[20];
    assign inter_3[17] = inter_2[17]^inter_2[21];
    assign inter_3[18] = inter_2[18]^inter_2[22];
    assign inter_3[19] = inter_2[19]^inter_2[23];
    assign inter_3[20] = inter_2[20];
    assign inter_3[21] = inter_2[21];
    assign inter_3[22] = inter_2[22];
    assign inter_3[23] = inter_2[23];
    assign inter_3[24] = inter_2[24]^inter_2[28];
    assign inter_3[25] = inter_2[25]^inter_2[29];
    assign inter_3[26] = inter_2[26]^inter_2[30];
    assign inter_3[27] = inter_2[27]^inter_2[31];
    assign inter_3[28] = inter_2[28];
    assign inter_3[29] = inter_2[29];
    assign inter_3[30] = inter_2[30];
    assign inter_3[31] = inter_2[31];
    assign inter_3[32] = inter_2[32]^inter_2[36];
    assign inter_3[33] = inter_2[33]^inter_2[37];
    assign inter_3[34] = inter_2[34]^inter_2[38];
    assign inter_3[35] = inter_2[35]^inter_2[39];
    assign inter_3[36] = inter_2[36];
    assign inter_3[37] = inter_2[37];
    assign inter_3[38] = inter_2[38];
    assign inter_3[39] = inter_2[39];
    assign inter_3[40] = inter_2[40]^inter_2[44];
    assign inter_3[41] = inter_2[41]^inter_2[45];
    assign inter_3[42] = inter_2[42]^inter_2[46];
    assign inter_3[43] = inter_2[43]^inter_2[47];
    assign inter_3[44] = inter_2[44];
    assign inter_3[45] = inter_2[45];
    assign inter_3[46] = inter_2[46];
    assign inter_3[47] = inter_2[47];
    assign inter_3[48] = inter_2[48]^inter_2[52];
    assign inter_3[49] = inter_2[49]^inter_2[53];
    assign inter_3[50] = inter_2[50]^inter_2[54];
    assign inter_3[51] = inter_2[51]^inter_2[55];
    assign inter_3[52] = inter_2[52];
    assign inter_3[53] = inter_2[53];
    assign inter_3[54] = inter_2[54];
    assign inter_3[55] = inter_2[55];
    assign inter_3[56] = inter_2[56]^inter_2[60];
    assign inter_3[57] = inter_2[57]^inter_2[61];
    assign inter_3[58] = inter_2[58]^inter_2[62];
    assign inter_3[59] = inter_2[59]^inter_2[63];
    assign inter_3[60] = inter_2[60];
    assign inter_3[61] = inter_2[61];
    assign inter_3[62] = inter_2[62];
    assign inter_3[63] = inter_2[63];
    assign inter_3[64] = inter_2[64]^inter_2[68];
    assign inter_3[65] = inter_2[65]^inter_2[69];
    assign inter_3[66] = inter_2[66]^inter_2[70];
    assign inter_3[67] = inter_2[67]^inter_2[71];
    assign inter_3[68] = inter_2[68];
    assign inter_3[69] = inter_2[69];
    assign inter_3[70] = inter_2[70];
    assign inter_3[71] = inter_2[71];
    assign inter_3[72] = inter_2[72]^inter_2[76];
    assign inter_3[73] = inter_2[73]^inter_2[77];
    assign inter_3[74] = inter_2[74]^inter_2[78];
    assign inter_3[75] = inter_2[75]^inter_2[79];
    assign inter_3[76] = inter_2[76];
    assign inter_3[77] = inter_2[77];
    assign inter_3[78] = inter_2[78];
    assign inter_3[79] = inter_2[79];
    assign inter_3[80] = inter_2[80]^inter_2[84];
    assign inter_3[81] = inter_2[81]^inter_2[85];
    assign inter_3[82] = inter_2[82]^inter_2[86];
    assign inter_3[83] = inter_2[83]^inter_2[87];
    assign inter_3[84] = inter_2[84];
    assign inter_3[85] = inter_2[85];
    assign inter_3[86] = inter_2[86];
    assign inter_3[87] = inter_2[87];
    assign inter_3[88] = inter_2[88]^inter_2[92];
    assign inter_3[89] = inter_2[89]^inter_2[93];
    assign inter_3[90] = inter_2[90]^inter_2[94];
    assign inter_3[91] = inter_2[91]^inter_2[95];
    assign inter_3[92] = inter_2[92];
    assign inter_3[93] = inter_2[93];
    assign inter_3[94] = inter_2[94];
    assign inter_3[95] = inter_2[95];
    assign inter_3[96] = inter_2[96]^inter_2[100];
    assign inter_3[97] = inter_2[97]^inter_2[101];
    assign inter_3[98] = inter_2[98]^inter_2[102];
    assign inter_3[99] = inter_2[99]^inter_2[103];
    assign inter_3[100] = inter_2[100];
    assign inter_3[101] = inter_2[101];
    assign inter_3[102] = inter_2[102];
    assign inter_3[103] = inter_2[103];
    assign inter_3[104] = inter_2[104]^inter_2[108];
    assign inter_3[105] = inter_2[105]^inter_2[109];
    assign inter_3[106] = inter_2[106]^inter_2[110];
    assign inter_3[107] = inter_2[107]^inter_2[111];
    assign inter_3[108] = inter_2[108];
    assign inter_3[109] = inter_2[109];
    assign inter_3[110] = inter_2[110];
    assign inter_3[111] = inter_2[111];
    assign inter_3[112] = inter_2[112]^inter_2[116];
    assign inter_3[113] = inter_2[113]^inter_2[117];
    assign inter_3[114] = inter_2[114]^inter_2[118];
    assign inter_3[115] = inter_2[115]^inter_2[119];
    assign inter_3[116] = inter_2[116];
    assign inter_3[117] = inter_2[117];
    assign inter_3[118] = inter_2[118];
    assign inter_3[119] = inter_2[119];
    assign inter_3[120] = inter_2[120]^inter_2[124];
    assign inter_3[121] = inter_2[121]^inter_2[125];
    assign inter_3[122] = inter_2[122]^inter_2[126];
    assign inter_3[123] = inter_2[123]^inter_2[127];
    assign inter_3[124] = inter_2[124];
    assign inter_3[125] = inter_2[125];
    assign inter_3[126] = inter_2[126];
    assign inter_3[127] = inter_2[127];
    assign inter_3[128] = inter_2[128]^inter_2[132];
    assign inter_3[129] = inter_2[129]^inter_2[133];
    assign inter_3[130] = inter_2[130]^inter_2[134];
    assign inter_3[131] = inter_2[131]^inter_2[135];
    assign inter_3[132] = inter_2[132];
    assign inter_3[133] = inter_2[133];
    assign inter_3[134] = inter_2[134];
    assign inter_3[135] = inter_2[135];
    assign inter_3[136] = inter_2[136]^inter_2[140];
    assign inter_3[137] = inter_2[137]^inter_2[141];
    assign inter_3[138] = inter_2[138]^inter_2[142];
    assign inter_3[139] = inter_2[139]^inter_2[143];
    assign inter_3[140] = inter_2[140];
    assign inter_3[141] = inter_2[141];
    assign inter_3[142] = inter_2[142];
    assign inter_3[143] = inter_2[143];
    assign inter_3[144] = inter_2[144]^inter_2[148];
    assign inter_3[145] = inter_2[145]^inter_2[149];
    assign inter_3[146] = inter_2[146]^inter_2[150];
    assign inter_3[147] = inter_2[147]^inter_2[151];
    assign inter_3[148] = inter_2[148];
    assign inter_3[149] = inter_2[149];
    assign inter_3[150] = inter_2[150];
    assign inter_3[151] = inter_2[151];
    assign inter_3[152] = inter_2[152]^inter_2[156];
    assign inter_3[153] = inter_2[153]^inter_2[157];
    assign inter_3[154] = inter_2[154]^inter_2[158];
    assign inter_3[155] = inter_2[155]^inter_2[159];
    assign inter_3[156] = inter_2[156];
    assign inter_3[157] = inter_2[157];
    assign inter_3[158] = inter_2[158];
    assign inter_3[159] = inter_2[159];
    assign inter_3[160] = inter_2[160]^inter_2[164];
    assign inter_3[161] = inter_2[161]^inter_2[165];
    assign inter_3[162] = inter_2[162]^inter_2[166];
    assign inter_3[163] = inter_2[163]^inter_2[167];
    assign inter_3[164] = inter_2[164];
    assign inter_3[165] = inter_2[165];
    assign inter_3[166] = inter_2[166];
    assign inter_3[167] = inter_2[167];
    assign inter_3[168] = inter_2[168]^inter_2[172];
    assign inter_3[169] = inter_2[169]^inter_2[173];
    assign inter_3[170] = inter_2[170]^inter_2[174];
    assign inter_3[171] = inter_2[171]^inter_2[175];
    assign inter_3[172] = inter_2[172];
    assign inter_3[173] = inter_2[173];
    assign inter_3[174] = inter_2[174];
    assign inter_3[175] = inter_2[175];
    assign inter_3[176] = inter_2[176]^inter_2[180];
    assign inter_3[177] = inter_2[177]^inter_2[181];
    assign inter_3[178] = inter_2[178]^inter_2[182];
    assign inter_3[179] = inter_2[179]^inter_2[183];
    assign inter_3[180] = inter_2[180];
    assign inter_3[181] = inter_2[181];
    assign inter_3[182] = inter_2[182];
    assign inter_3[183] = inter_2[183];
    assign inter_3[184] = inter_2[184]^inter_2[188];
    assign inter_3[185] = inter_2[185]^inter_2[189];
    assign inter_3[186] = inter_2[186]^inter_2[190];
    assign inter_3[187] = inter_2[187]^inter_2[191];
    assign inter_3[188] = inter_2[188];
    assign inter_3[189] = inter_2[189];
    assign inter_3[190] = inter_2[190];
    assign inter_3[191] = inter_2[191];
    assign inter_3[192] = inter_2[192]^inter_2[196];
    assign inter_3[193] = inter_2[193]^inter_2[197];
    assign inter_3[194] = inter_2[194]^inter_2[198];
    assign inter_3[195] = inter_2[195]^inter_2[199];
    assign inter_3[196] = inter_2[196];
    assign inter_3[197] = inter_2[197];
    assign inter_3[198] = inter_2[198];
    assign inter_3[199] = inter_2[199];
    assign inter_3[200] = inter_2[200]^inter_2[204];
    assign inter_3[201] = inter_2[201]^inter_2[205];
    assign inter_3[202] = inter_2[202]^inter_2[206];
    assign inter_3[203] = inter_2[203]^inter_2[207];
    assign inter_3[204] = inter_2[204];
    assign inter_3[205] = inter_2[205];
    assign inter_3[206] = inter_2[206];
    assign inter_3[207] = inter_2[207];
    assign inter_3[208] = inter_2[208]^inter_2[212];
    assign inter_3[209] = inter_2[209]^inter_2[213];
    assign inter_3[210] = inter_2[210]^inter_2[214];
    assign inter_3[211] = inter_2[211]^inter_2[215];
    assign inter_3[212] = inter_2[212];
    assign inter_3[213] = inter_2[213];
    assign inter_3[214] = inter_2[214];
    assign inter_3[215] = inter_2[215];
    assign inter_3[216] = inter_2[216]^inter_2[220];
    assign inter_3[217] = inter_2[217]^inter_2[221];
    assign inter_3[218] = inter_2[218]^inter_2[222];
    assign inter_3[219] = inter_2[219]^inter_2[223];
    assign inter_3[220] = inter_2[220];
    assign inter_3[221] = inter_2[221];
    assign inter_3[222] = inter_2[222];
    assign inter_3[223] = inter_2[223];
    assign inter_3[224] = inter_2[224]^inter_2[228];
    assign inter_3[225] = inter_2[225]^inter_2[229];
    assign inter_3[226] = inter_2[226]^inter_2[230];
    assign inter_3[227] = inter_2[227]^inter_2[231];
    assign inter_3[228] = inter_2[228];
    assign inter_3[229] = inter_2[229];
    assign inter_3[230] = inter_2[230];
    assign inter_3[231] = inter_2[231];
    assign inter_3[232] = inter_2[232]^inter_2[236];
    assign inter_3[233] = inter_2[233]^inter_2[237];
    assign inter_3[234] = inter_2[234]^inter_2[238];
    assign inter_3[235] = inter_2[235]^inter_2[239];
    assign inter_3[236] = inter_2[236];
    assign inter_3[237] = inter_2[237];
    assign inter_3[238] = inter_2[238];
    assign inter_3[239] = inter_2[239];
    assign inter_3[240] = inter_2[240]^inter_2[244];
    assign inter_3[241] = inter_2[241]^inter_2[245];
    assign inter_3[242] = inter_2[242]^inter_2[246];
    assign inter_3[243] = inter_2[243]^inter_2[247];
    assign inter_3[244] = inter_2[244];
    assign inter_3[245] = inter_2[245];
    assign inter_3[246] = inter_2[246];
    assign inter_3[247] = inter_2[247];
    assign inter_3[248] = inter_2[248]^inter_2[252];
    assign inter_3[249] = inter_2[249]^inter_2[253];
    assign inter_3[250] = inter_2[250]^inter_2[254];
    assign inter_3[251] = inter_2[251]^inter_2[255];
    assign inter_3[252] = inter_2[252];
    assign inter_3[253] = inter_2[253];
    assign inter_3[254] = inter_2[254];
    assign inter_3[255] = inter_2[255];
    assign inter_3[256] = inter_2[256]^inter_2[260];
    assign inter_3[257] = inter_2[257]^inter_2[261];
    assign inter_3[258] = inter_2[258]^inter_2[262];
    assign inter_3[259] = inter_2[259]^inter_2[263];
    assign inter_3[260] = inter_2[260];
    assign inter_3[261] = inter_2[261];
    assign inter_3[262] = inter_2[262];
    assign inter_3[263] = inter_2[263];
    assign inter_3[264] = inter_2[264]^inter_2[268];
    assign inter_3[265] = inter_2[265]^inter_2[269];
    assign inter_3[266] = inter_2[266]^inter_2[270];
    assign inter_3[267] = inter_2[267]^inter_2[271];
    assign inter_3[268] = inter_2[268];
    assign inter_3[269] = inter_2[269];
    assign inter_3[270] = inter_2[270];
    assign inter_3[271] = inter_2[271];
    assign inter_3[272] = inter_2[272]^inter_2[276];
    assign inter_3[273] = inter_2[273]^inter_2[277];
    assign inter_3[274] = inter_2[274]^inter_2[278];
    assign inter_3[275] = inter_2[275]^inter_2[279];
    assign inter_3[276] = inter_2[276];
    assign inter_3[277] = inter_2[277];
    assign inter_3[278] = inter_2[278];
    assign inter_3[279] = inter_2[279];
    assign inter_3[280] = inter_2[280]^inter_2[284];
    assign inter_3[281] = inter_2[281]^inter_2[285];
    assign inter_3[282] = inter_2[282]^inter_2[286];
    assign inter_3[283] = inter_2[283]^inter_2[287];
    assign inter_3[284] = inter_2[284];
    assign inter_3[285] = inter_2[285];
    assign inter_3[286] = inter_2[286];
    assign inter_3[287] = inter_2[287];
    assign inter_3[288] = inter_2[288]^inter_2[292];
    assign inter_3[289] = inter_2[289]^inter_2[293];
    assign inter_3[290] = inter_2[290]^inter_2[294];
    assign inter_3[291] = inter_2[291]^inter_2[295];
    assign inter_3[292] = inter_2[292];
    assign inter_3[293] = inter_2[293];
    assign inter_3[294] = inter_2[294];
    assign inter_3[295] = inter_2[295];
    assign inter_3[296] = inter_2[296]^inter_2[300];
    assign inter_3[297] = inter_2[297]^inter_2[301];
    assign inter_3[298] = inter_2[298]^inter_2[302];
    assign inter_3[299] = inter_2[299]^inter_2[303];
    assign inter_3[300] = inter_2[300];
    assign inter_3[301] = inter_2[301];
    assign inter_3[302] = inter_2[302];
    assign inter_3[303] = inter_2[303];
    assign inter_3[304] = inter_2[304]^inter_2[308];
    assign inter_3[305] = inter_2[305]^inter_2[309];
    assign inter_3[306] = inter_2[306]^inter_2[310];
    assign inter_3[307] = inter_2[307]^inter_2[311];
    assign inter_3[308] = inter_2[308];
    assign inter_3[309] = inter_2[309];
    assign inter_3[310] = inter_2[310];
    assign inter_3[311] = inter_2[311];
    assign inter_3[312] = inter_2[312]^inter_2[316];
    assign inter_3[313] = inter_2[313]^inter_2[317];
    assign inter_3[314] = inter_2[314]^inter_2[318];
    assign inter_3[315] = inter_2[315]^inter_2[319];
    assign inter_3[316] = inter_2[316];
    assign inter_3[317] = inter_2[317];
    assign inter_3[318] = inter_2[318];
    assign inter_3[319] = inter_2[319];
    assign inter_3[320] = inter_2[320]^inter_2[324];
    assign inter_3[321] = inter_2[321]^inter_2[325];
    assign inter_3[322] = inter_2[322]^inter_2[326];
    assign inter_3[323] = inter_2[323]^inter_2[327];
    assign inter_3[324] = inter_2[324];
    assign inter_3[325] = inter_2[325];
    assign inter_3[326] = inter_2[326];
    assign inter_3[327] = inter_2[327];
    assign inter_3[328] = inter_2[328]^inter_2[332];
    assign inter_3[329] = inter_2[329]^inter_2[333];
    assign inter_3[330] = inter_2[330]^inter_2[334];
    assign inter_3[331] = inter_2[331]^inter_2[335];
    assign inter_3[332] = inter_2[332];
    assign inter_3[333] = inter_2[333];
    assign inter_3[334] = inter_2[334];
    assign inter_3[335] = inter_2[335];
    assign inter_3[336] = inter_2[336]^inter_2[340];
    assign inter_3[337] = inter_2[337]^inter_2[341];
    assign inter_3[338] = inter_2[338]^inter_2[342];
    assign inter_3[339] = inter_2[339]^inter_2[343];
    assign inter_3[340] = inter_2[340];
    assign inter_3[341] = inter_2[341];
    assign inter_3[342] = inter_2[342];
    assign inter_3[343] = inter_2[343];
    assign inter_3[344] = inter_2[344]^inter_2[348];
    assign inter_3[345] = inter_2[345]^inter_2[349];
    assign inter_3[346] = inter_2[346]^inter_2[350];
    assign inter_3[347] = inter_2[347]^inter_2[351];
    assign inter_3[348] = inter_2[348];
    assign inter_3[349] = inter_2[349];
    assign inter_3[350] = inter_2[350];
    assign inter_3[351] = inter_2[351];
    assign inter_3[352] = inter_2[352]^inter_2[356];
    assign inter_3[353] = inter_2[353]^inter_2[357];
    assign inter_3[354] = inter_2[354]^inter_2[358];
    assign inter_3[355] = inter_2[355]^inter_2[359];
    assign inter_3[356] = inter_2[356];
    assign inter_3[357] = inter_2[357];
    assign inter_3[358] = inter_2[358];
    assign inter_3[359] = inter_2[359];
    assign inter_3[360] = inter_2[360]^inter_2[364];
    assign inter_3[361] = inter_2[361]^inter_2[365];
    assign inter_3[362] = inter_2[362]^inter_2[366];
    assign inter_3[363] = inter_2[363]^inter_2[367];
    assign inter_3[364] = inter_2[364];
    assign inter_3[365] = inter_2[365];
    assign inter_3[366] = inter_2[366];
    assign inter_3[367] = inter_2[367];
    assign inter_3[368] = inter_2[368]^inter_2[372];
    assign inter_3[369] = inter_2[369]^inter_2[373];
    assign inter_3[370] = inter_2[370]^inter_2[374];
    assign inter_3[371] = inter_2[371]^inter_2[375];
    assign inter_3[372] = inter_2[372];
    assign inter_3[373] = inter_2[373];
    assign inter_3[374] = inter_2[374];
    assign inter_3[375] = inter_2[375];
    assign inter_3[376] = inter_2[376]^inter_2[380];
    assign inter_3[377] = inter_2[377]^inter_2[381];
    assign inter_3[378] = inter_2[378]^inter_2[382];
    assign inter_3[379] = inter_2[379]^inter_2[383];
    assign inter_3[380] = inter_2[380];
    assign inter_3[381] = inter_2[381];
    assign inter_3[382] = inter_2[382];
    assign inter_3[383] = inter_2[383];
    assign inter_3[384] = inter_2[384]^inter_2[388];
    assign inter_3[385] = inter_2[385]^inter_2[389];
    assign inter_3[386] = inter_2[386]^inter_2[390];
    assign inter_3[387] = inter_2[387]^inter_2[391];
    assign inter_3[388] = inter_2[388];
    assign inter_3[389] = inter_2[389];
    assign inter_3[390] = inter_2[390];
    assign inter_3[391] = inter_2[391];
    assign inter_3[392] = inter_2[392]^inter_2[396];
    assign inter_3[393] = inter_2[393]^inter_2[397];
    assign inter_3[394] = inter_2[394]^inter_2[398];
    assign inter_3[395] = inter_2[395]^inter_2[399];
    assign inter_3[396] = inter_2[396];
    assign inter_3[397] = inter_2[397];
    assign inter_3[398] = inter_2[398];
    assign inter_3[399] = inter_2[399];
    assign inter_3[400] = inter_2[400]^inter_2[404];
    assign inter_3[401] = inter_2[401]^inter_2[405];
    assign inter_3[402] = inter_2[402]^inter_2[406];
    assign inter_3[403] = inter_2[403]^inter_2[407];
    assign inter_3[404] = inter_2[404];
    assign inter_3[405] = inter_2[405];
    assign inter_3[406] = inter_2[406];
    assign inter_3[407] = inter_2[407];
    assign inter_3[408] = inter_2[408]^inter_2[412];
    assign inter_3[409] = inter_2[409]^inter_2[413];
    assign inter_3[410] = inter_2[410]^inter_2[414];
    assign inter_3[411] = inter_2[411]^inter_2[415];
    assign inter_3[412] = inter_2[412];
    assign inter_3[413] = inter_2[413];
    assign inter_3[414] = inter_2[414];
    assign inter_3[415] = inter_2[415];
    assign inter_3[416] = inter_2[416]^inter_2[420];
    assign inter_3[417] = inter_2[417]^inter_2[421];
    assign inter_3[418] = inter_2[418]^inter_2[422];
    assign inter_3[419] = inter_2[419]^inter_2[423];
    assign inter_3[420] = inter_2[420];
    assign inter_3[421] = inter_2[421];
    assign inter_3[422] = inter_2[422];
    assign inter_3[423] = inter_2[423];
    assign inter_3[424] = inter_2[424]^inter_2[428];
    assign inter_3[425] = inter_2[425]^inter_2[429];
    assign inter_3[426] = inter_2[426]^inter_2[430];
    assign inter_3[427] = inter_2[427]^inter_2[431];
    assign inter_3[428] = inter_2[428];
    assign inter_3[429] = inter_2[429];
    assign inter_3[430] = inter_2[430];
    assign inter_3[431] = inter_2[431];
    assign inter_3[432] = inter_2[432]^inter_2[436];
    assign inter_3[433] = inter_2[433]^inter_2[437];
    assign inter_3[434] = inter_2[434]^inter_2[438];
    assign inter_3[435] = inter_2[435]^inter_2[439];
    assign inter_3[436] = inter_2[436];
    assign inter_3[437] = inter_2[437];
    assign inter_3[438] = inter_2[438];
    assign inter_3[439] = inter_2[439];
    assign inter_3[440] = inter_2[440]^inter_2[444];
    assign inter_3[441] = inter_2[441]^inter_2[445];
    assign inter_3[442] = inter_2[442]^inter_2[446];
    assign inter_3[443] = inter_2[443]^inter_2[447];
    assign inter_3[444] = inter_2[444];
    assign inter_3[445] = inter_2[445];
    assign inter_3[446] = inter_2[446];
    assign inter_3[447] = inter_2[447];
    assign inter_3[448] = inter_2[448]^inter_2[452];
    assign inter_3[449] = inter_2[449]^inter_2[453];
    assign inter_3[450] = inter_2[450]^inter_2[454];
    assign inter_3[451] = inter_2[451]^inter_2[455];
    assign inter_3[452] = inter_2[452];
    assign inter_3[453] = inter_2[453];
    assign inter_3[454] = inter_2[454];
    assign inter_3[455] = inter_2[455];
    assign inter_3[456] = inter_2[456]^inter_2[460];
    assign inter_3[457] = inter_2[457]^inter_2[461];
    assign inter_3[458] = inter_2[458]^inter_2[462];
    assign inter_3[459] = inter_2[459]^inter_2[463];
    assign inter_3[460] = inter_2[460];
    assign inter_3[461] = inter_2[461];
    assign inter_3[462] = inter_2[462];
    assign inter_3[463] = inter_2[463];
    assign inter_3[464] = inter_2[464]^inter_2[468];
    assign inter_3[465] = inter_2[465]^inter_2[469];
    assign inter_3[466] = inter_2[466]^inter_2[470];
    assign inter_3[467] = inter_2[467]^inter_2[471];
    assign inter_3[468] = inter_2[468];
    assign inter_3[469] = inter_2[469];
    assign inter_3[470] = inter_2[470];
    assign inter_3[471] = inter_2[471];
    assign inter_3[472] = inter_2[472]^inter_2[476];
    assign inter_3[473] = inter_2[473]^inter_2[477];
    assign inter_3[474] = inter_2[474]^inter_2[478];
    assign inter_3[475] = inter_2[475]^inter_2[479];
    assign inter_3[476] = inter_2[476];
    assign inter_3[477] = inter_2[477];
    assign inter_3[478] = inter_2[478];
    assign inter_3[479] = inter_2[479];
    assign inter_3[480] = inter_2[480]^inter_2[484];
    assign inter_3[481] = inter_2[481]^inter_2[485];
    assign inter_3[482] = inter_2[482]^inter_2[486];
    assign inter_3[483] = inter_2[483]^inter_2[487];
    assign inter_3[484] = inter_2[484];
    assign inter_3[485] = inter_2[485];
    assign inter_3[486] = inter_2[486];
    assign inter_3[487] = inter_2[487];
    assign inter_3[488] = inter_2[488]^inter_2[492];
    assign inter_3[489] = inter_2[489]^inter_2[493];
    assign inter_3[490] = inter_2[490]^inter_2[494];
    assign inter_3[491] = inter_2[491]^inter_2[495];
    assign inter_3[492] = inter_2[492];
    assign inter_3[493] = inter_2[493];
    assign inter_3[494] = inter_2[494];
    assign inter_3[495] = inter_2[495];
    assign inter_3[496] = inter_2[496]^inter_2[500];
    assign inter_3[497] = inter_2[497]^inter_2[501];
    assign inter_3[498] = inter_2[498]^inter_2[502];
    assign inter_3[499] = inter_2[499]^inter_2[503];
    assign inter_3[500] = inter_2[500];
    assign inter_3[501] = inter_2[501];
    assign inter_3[502] = inter_2[502];
    assign inter_3[503] = inter_2[503];
    assign inter_3[504] = inter_2[504]^inter_2[508];
    assign inter_3[505] = inter_2[505]^inter_2[509];
    assign inter_3[506] = inter_2[506]^inter_2[510];
    assign inter_3[507] = inter_2[507]^inter_2[511];
    assign inter_3[508] = inter_2[508];
    assign inter_3[509] = inter_2[509];
    assign inter_3[510] = inter_2[510];
    assign inter_3[511] = inter_2[511];
    assign inter_3[512] = inter_2[512]^inter_2[516];
    assign inter_3[513] = inter_2[513]^inter_2[517];
    assign inter_3[514] = inter_2[514]^inter_2[518];
    assign inter_3[515] = inter_2[515]^inter_2[519];
    assign inter_3[516] = inter_2[516];
    assign inter_3[517] = inter_2[517];
    assign inter_3[518] = inter_2[518];
    assign inter_3[519] = inter_2[519];
    assign inter_3[520] = inter_2[520]^inter_2[524];
    assign inter_3[521] = inter_2[521]^inter_2[525];
    assign inter_3[522] = inter_2[522]^inter_2[526];
    assign inter_3[523] = inter_2[523]^inter_2[527];
    assign inter_3[524] = inter_2[524];
    assign inter_3[525] = inter_2[525];
    assign inter_3[526] = inter_2[526];
    assign inter_3[527] = inter_2[527];
    assign inter_3[528] = inter_2[528]^inter_2[532];
    assign inter_3[529] = inter_2[529]^inter_2[533];
    assign inter_3[530] = inter_2[530]^inter_2[534];
    assign inter_3[531] = inter_2[531]^inter_2[535];
    assign inter_3[532] = inter_2[532];
    assign inter_3[533] = inter_2[533];
    assign inter_3[534] = inter_2[534];
    assign inter_3[535] = inter_2[535];
    assign inter_3[536] = inter_2[536]^inter_2[540];
    assign inter_3[537] = inter_2[537]^inter_2[541];
    assign inter_3[538] = inter_2[538]^inter_2[542];
    assign inter_3[539] = inter_2[539]^inter_2[543];
    assign inter_3[540] = inter_2[540];
    assign inter_3[541] = inter_2[541];
    assign inter_3[542] = inter_2[542];
    assign inter_3[543] = inter_2[543];
    assign inter_3[544] = inter_2[544]^inter_2[548];
    assign inter_3[545] = inter_2[545]^inter_2[549];
    assign inter_3[546] = inter_2[546]^inter_2[550];
    assign inter_3[547] = inter_2[547]^inter_2[551];
    assign inter_3[548] = inter_2[548];
    assign inter_3[549] = inter_2[549];
    assign inter_3[550] = inter_2[550];
    assign inter_3[551] = inter_2[551];
    assign inter_3[552] = inter_2[552]^inter_2[556];
    assign inter_3[553] = inter_2[553]^inter_2[557];
    assign inter_3[554] = inter_2[554]^inter_2[558];
    assign inter_3[555] = inter_2[555]^inter_2[559];
    assign inter_3[556] = inter_2[556];
    assign inter_3[557] = inter_2[557];
    assign inter_3[558] = inter_2[558];
    assign inter_3[559] = inter_2[559];
    assign inter_3[560] = inter_2[560]^inter_2[564];
    assign inter_3[561] = inter_2[561]^inter_2[565];
    assign inter_3[562] = inter_2[562]^inter_2[566];
    assign inter_3[563] = inter_2[563]^inter_2[567];
    assign inter_3[564] = inter_2[564];
    assign inter_3[565] = inter_2[565];
    assign inter_3[566] = inter_2[566];
    assign inter_3[567] = inter_2[567];
    assign inter_3[568] = inter_2[568]^inter_2[572];
    assign inter_3[569] = inter_2[569]^inter_2[573];
    assign inter_3[570] = inter_2[570]^inter_2[574];
    assign inter_3[571] = inter_2[571]^inter_2[575];
    assign inter_3[572] = inter_2[572];
    assign inter_3[573] = inter_2[573];
    assign inter_3[574] = inter_2[574];
    assign inter_3[575] = inter_2[575];
    assign inter_3[576] = inter_2[576]^inter_2[580];
    assign inter_3[577] = inter_2[577]^inter_2[581];
    assign inter_3[578] = inter_2[578]^inter_2[582];
    assign inter_3[579] = inter_2[579]^inter_2[583];
    assign inter_3[580] = inter_2[580];
    assign inter_3[581] = inter_2[581];
    assign inter_3[582] = inter_2[582];
    assign inter_3[583] = inter_2[583];
    assign inter_3[584] = inter_2[584]^inter_2[588];
    assign inter_3[585] = inter_2[585]^inter_2[589];
    assign inter_3[586] = inter_2[586]^inter_2[590];
    assign inter_3[587] = inter_2[587]^inter_2[591];
    assign inter_3[588] = inter_2[588];
    assign inter_3[589] = inter_2[589];
    assign inter_3[590] = inter_2[590];
    assign inter_3[591] = inter_2[591];
    assign inter_3[592] = inter_2[592]^inter_2[596];
    assign inter_3[593] = inter_2[593]^inter_2[597];
    assign inter_3[594] = inter_2[594]^inter_2[598];
    assign inter_3[595] = inter_2[595]^inter_2[599];
    assign inter_3[596] = inter_2[596];
    assign inter_3[597] = inter_2[597];
    assign inter_3[598] = inter_2[598];
    assign inter_3[599] = inter_2[599];
    assign inter_3[600] = inter_2[600]^inter_2[604];
    assign inter_3[601] = inter_2[601]^inter_2[605];
    assign inter_3[602] = inter_2[602]^inter_2[606];
    assign inter_3[603] = inter_2[603]^inter_2[607];
    assign inter_3[604] = inter_2[604];
    assign inter_3[605] = inter_2[605];
    assign inter_3[606] = inter_2[606];
    assign inter_3[607] = inter_2[607];
    assign inter_3[608] = inter_2[608]^inter_2[612];
    assign inter_3[609] = inter_2[609]^inter_2[613];
    assign inter_3[610] = inter_2[610]^inter_2[614];
    assign inter_3[611] = inter_2[611]^inter_2[615];
    assign inter_3[612] = inter_2[612];
    assign inter_3[613] = inter_2[613];
    assign inter_3[614] = inter_2[614];
    assign inter_3[615] = inter_2[615];
    assign inter_3[616] = inter_2[616]^inter_2[620];
    assign inter_3[617] = inter_2[617]^inter_2[621];
    assign inter_3[618] = inter_2[618]^inter_2[622];
    assign inter_3[619] = inter_2[619]^inter_2[623];
    assign inter_3[620] = inter_2[620];
    assign inter_3[621] = inter_2[621];
    assign inter_3[622] = inter_2[622];
    assign inter_3[623] = inter_2[623];
    assign inter_3[624] = inter_2[624]^inter_2[628];
    assign inter_3[625] = inter_2[625]^inter_2[629];
    assign inter_3[626] = inter_2[626]^inter_2[630];
    assign inter_3[627] = inter_2[627]^inter_2[631];
    assign inter_3[628] = inter_2[628];
    assign inter_3[629] = inter_2[629];
    assign inter_3[630] = inter_2[630];
    assign inter_3[631] = inter_2[631];
    assign inter_3[632] = inter_2[632]^inter_2[636];
    assign inter_3[633] = inter_2[633]^inter_2[637];
    assign inter_3[634] = inter_2[634]^inter_2[638];
    assign inter_3[635] = inter_2[635]^inter_2[639];
    assign inter_3[636] = inter_2[636];
    assign inter_3[637] = inter_2[637];
    assign inter_3[638] = inter_2[638];
    assign inter_3[639] = inter_2[639];
    assign inter_3[640] = inter_2[640]^inter_2[644];
    assign inter_3[641] = inter_2[641]^inter_2[645];
    assign inter_3[642] = inter_2[642]^inter_2[646];
    assign inter_3[643] = inter_2[643]^inter_2[647];
    assign inter_3[644] = inter_2[644];
    assign inter_3[645] = inter_2[645];
    assign inter_3[646] = inter_2[646];
    assign inter_3[647] = inter_2[647];
    assign inter_3[648] = inter_2[648]^inter_2[652];
    assign inter_3[649] = inter_2[649]^inter_2[653];
    assign inter_3[650] = inter_2[650]^inter_2[654];
    assign inter_3[651] = inter_2[651]^inter_2[655];
    assign inter_3[652] = inter_2[652];
    assign inter_3[653] = inter_2[653];
    assign inter_3[654] = inter_2[654];
    assign inter_3[655] = inter_2[655];
    assign inter_3[656] = inter_2[656]^inter_2[660];
    assign inter_3[657] = inter_2[657]^inter_2[661];
    assign inter_3[658] = inter_2[658]^inter_2[662];
    assign inter_3[659] = inter_2[659]^inter_2[663];
    assign inter_3[660] = inter_2[660];
    assign inter_3[661] = inter_2[661];
    assign inter_3[662] = inter_2[662];
    assign inter_3[663] = inter_2[663];
    assign inter_3[664] = inter_2[664]^inter_2[668];
    assign inter_3[665] = inter_2[665]^inter_2[669];
    assign inter_3[666] = inter_2[666]^inter_2[670];
    assign inter_3[667] = inter_2[667]^inter_2[671];
    assign inter_3[668] = inter_2[668];
    assign inter_3[669] = inter_2[669];
    assign inter_3[670] = inter_2[670];
    assign inter_3[671] = inter_2[671];
    assign inter_3[672] = inter_2[672]^inter_2[676];
    assign inter_3[673] = inter_2[673]^inter_2[677];
    assign inter_3[674] = inter_2[674]^inter_2[678];
    assign inter_3[675] = inter_2[675]^inter_2[679];
    assign inter_3[676] = inter_2[676];
    assign inter_3[677] = inter_2[677];
    assign inter_3[678] = inter_2[678];
    assign inter_3[679] = inter_2[679];
    assign inter_3[680] = inter_2[680]^inter_2[684];
    assign inter_3[681] = inter_2[681]^inter_2[685];
    assign inter_3[682] = inter_2[682]^inter_2[686];
    assign inter_3[683] = inter_2[683]^inter_2[687];
    assign inter_3[684] = inter_2[684];
    assign inter_3[685] = inter_2[685];
    assign inter_3[686] = inter_2[686];
    assign inter_3[687] = inter_2[687];
    assign inter_3[688] = inter_2[688]^inter_2[692];
    assign inter_3[689] = inter_2[689]^inter_2[693];
    assign inter_3[690] = inter_2[690]^inter_2[694];
    assign inter_3[691] = inter_2[691]^inter_2[695];
    assign inter_3[692] = inter_2[692];
    assign inter_3[693] = inter_2[693];
    assign inter_3[694] = inter_2[694];
    assign inter_3[695] = inter_2[695];
    assign inter_3[696] = inter_2[696]^inter_2[700];
    assign inter_3[697] = inter_2[697]^inter_2[701];
    assign inter_3[698] = inter_2[698]^inter_2[702];
    assign inter_3[699] = inter_2[699]^inter_2[703];
    assign inter_3[700] = inter_2[700];
    assign inter_3[701] = inter_2[701];
    assign inter_3[702] = inter_2[702];
    assign inter_3[703] = inter_2[703];
    assign inter_3[704] = inter_2[704]^inter_2[708];
    assign inter_3[705] = inter_2[705]^inter_2[709];
    assign inter_3[706] = inter_2[706]^inter_2[710];
    assign inter_3[707] = inter_2[707]^inter_2[711];
    assign inter_3[708] = inter_2[708];
    assign inter_3[709] = inter_2[709];
    assign inter_3[710] = inter_2[710];
    assign inter_3[711] = inter_2[711];
    assign inter_3[712] = inter_2[712]^inter_2[716];
    assign inter_3[713] = inter_2[713]^inter_2[717];
    assign inter_3[714] = inter_2[714]^inter_2[718];
    assign inter_3[715] = inter_2[715]^inter_2[719];
    assign inter_3[716] = inter_2[716];
    assign inter_3[717] = inter_2[717];
    assign inter_3[718] = inter_2[718];
    assign inter_3[719] = inter_2[719];
    assign inter_3[720] = inter_2[720]^inter_2[724];
    assign inter_3[721] = inter_2[721]^inter_2[725];
    assign inter_3[722] = inter_2[722]^inter_2[726];
    assign inter_3[723] = inter_2[723]^inter_2[727];
    assign inter_3[724] = inter_2[724];
    assign inter_3[725] = inter_2[725];
    assign inter_3[726] = inter_2[726];
    assign inter_3[727] = inter_2[727];
    assign inter_3[728] = inter_2[728]^inter_2[732];
    assign inter_3[729] = inter_2[729]^inter_2[733];
    assign inter_3[730] = inter_2[730]^inter_2[734];
    assign inter_3[731] = inter_2[731]^inter_2[735];
    assign inter_3[732] = inter_2[732];
    assign inter_3[733] = inter_2[733];
    assign inter_3[734] = inter_2[734];
    assign inter_3[735] = inter_2[735];
    assign inter_3[736] = inter_2[736]^inter_2[740];
    assign inter_3[737] = inter_2[737]^inter_2[741];
    assign inter_3[738] = inter_2[738]^inter_2[742];
    assign inter_3[739] = inter_2[739]^inter_2[743];
    assign inter_3[740] = inter_2[740];
    assign inter_3[741] = inter_2[741];
    assign inter_3[742] = inter_2[742];
    assign inter_3[743] = inter_2[743];
    assign inter_3[744] = inter_2[744]^inter_2[748];
    assign inter_3[745] = inter_2[745]^inter_2[749];
    assign inter_3[746] = inter_2[746]^inter_2[750];
    assign inter_3[747] = inter_2[747]^inter_2[751];
    assign inter_3[748] = inter_2[748];
    assign inter_3[749] = inter_2[749];
    assign inter_3[750] = inter_2[750];
    assign inter_3[751] = inter_2[751];
    assign inter_3[752] = inter_2[752]^inter_2[756];
    assign inter_3[753] = inter_2[753]^inter_2[757];
    assign inter_3[754] = inter_2[754]^inter_2[758];
    assign inter_3[755] = inter_2[755]^inter_2[759];
    assign inter_3[756] = inter_2[756];
    assign inter_3[757] = inter_2[757];
    assign inter_3[758] = inter_2[758];
    assign inter_3[759] = inter_2[759];
    assign inter_3[760] = inter_2[760]^inter_2[764];
    assign inter_3[761] = inter_2[761]^inter_2[765];
    assign inter_3[762] = inter_2[762]^inter_2[766];
    assign inter_3[763] = inter_2[763]^inter_2[767];
    assign inter_3[764] = inter_2[764];
    assign inter_3[765] = inter_2[765];
    assign inter_3[766] = inter_2[766];
    assign inter_3[767] = inter_2[767];
    assign inter_3[768] = inter_2[768]^inter_2[772];
    assign inter_3[769] = inter_2[769]^inter_2[773];
    assign inter_3[770] = inter_2[770]^inter_2[774];
    assign inter_3[771] = inter_2[771]^inter_2[775];
    assign inter_3[772] = inter_2[772];
    assign inter_3[773] = inter_2[773];
    assign inter_3[774] = inter_2[774];
    assign inter_3[775] = inter_2[775];
    assign inter_3[776] = inter_2[776]^inter_2[780];
    assign inter_3[777] = inter_2[777]^inter_2[781];
    assign inter_3[778] = inter_2[778]^inter_2[782];
    assign inter_3[779] = inter_2[779]^inter_2[783];
    assign inter_3[780] = inter_2[780];
    assign inter_3[781] = inter_2[781];
    assign inter_3[782] = inter_2[782];
    assign inter_3[783] = inter_2[783];
    assign inter_3[784] = inter_2[784]^inter_2[788];
    assign inter_3[785] = inter_2[785]^inter_2[789];
    assign inter_3[786] = inter_2[786]^inter_2[790];
    assign inter_3[787] = inter_2[787]^inter_2[791];
    assign inter_3[788] = inter_2[788];
    assign inter_3[789] = inter_2[789];
    assign inter_3[790] = inter_2[790];
    assign inter_3[791] = inter_2[791];
    assign inter_3[792] = inter_2[792]^inter_2[796];
    assign inter_3[793] = inter_2[793]^inter_2[797];
    assign inter_3[794] = inter_2[794]^inter_2[798];
    assign inter_3[795] = inter_2[795]^inter_2[799];
    assign inter_3[796] = inter_2[796];
    assign inter_3[797] = inter_2[797];
    assign inter_3[798] = inter_2[798];
    assign inter_3[799] = inter_2[799];
    assign inter_3[800] = inter_2[800]^inter_2[804];
    assign inter_3[801] = inter_2[801]^inter_2[805];
    assign inter_3[802] = inter_2[802]^inter_2[806];
    assign inter_3[803] = inter_2[803]^inter_2[807];
    assign inter_3[804] = inter_2[804];
    assign inter_3[805] = inter_2[805];
    assign inter_3[806] = inter_2[806];
    assign inter_3[807] = inter_2[807];
    assign inter_3[808] = inter_2[808]^inter_2[812];
    assign inter_3[809] = inter_2[809]^inter_2[813];
    assign inter_3[810] = inter_2[810]^inter_2[814];
    assign inter_3[811] = inter_2[811]^inter_2[815];
    assign inter_3[812] = inter_2[812];
    assign inter_3[813] = inter_2[813];
    assign inter_3[814] = inter_2[814];
    assign inter_3[815] = inter_2[815];
    assign inter_3[816] = inter_2[816]^inter_2[820];
    assign inter_3[817] = inter_2[817]^inter_2[821];
    assign inter_3[818] = inter_2[818]^inter_2[822];
    assign inter_3[819] = inter_2[819]^inter_2[823];
    assign inter_3[820] = inter_2[820];
    assign inter_3[821] = inter_2[821];
    assign inter_3[822] = inter_2[822];
    assign inter_3[823] = inter_2[823];
    assign inter_3[824] = inter_2[824]^inter_2[828];
    assign inter_3[825] = inter_2[825]^inter_2[829];
    assign inter_3[826] = inter_2[826]^inter_2[830];
    assign inter_3[827] = inter_2[827]^inter_2[831];
    assign inter_3[828] = inter_2[828];
    assign inter_3[829] = inter_2[829];
    assign inter_3[830] = inter_2[830];
    assign inter_3[831] = inter_2[831];
    assign inter_3[832] = inter_2[832]^inter_2[836];
    assign inter_3[833] = inter_2[833]^inter_2[837];
    assign inter_3[834] = inter_2[834]^inter_2[838];
    assign inter_3[835] = inter_2[835]^inter_2[839];
    assign inter_3[836] = inter_2[836];
    assign inter_3[837] = inter_2[837];
    assign inter_3[838] = inter_2[838];
    assign inter_3[839] = inter_2[839];
    assign inter_3[840] = inter_2[840]^inter_2[844];
    assign inter_3[841] = inter_2[841]^inter_2[845];
    assign inter_3[842] = inter_2[842]^inter_2[846];
    assign inter_3[843] = inter_2[843]^inter_2[847];
    assign inter_3[844] = inter_2[844];
    assign inter_3[845] = inter_2[845];
    assign inter_3[846] = inter_2[846];
    assign inter_3[847] = inter_2[847];
    assign inter_3[848] = inter_2[848]^inter_2[852];
    assign inter_3[849] = inter_2[849]^inter_2[853];
    assign inter_3[850] = inter_2[850]^inter_2[854];
    assign inter_3[851] = inter_2[851]^inter_2[855];
    assign inter_3[852] = inter_2[852];
    assign inter_3[853] = inter_2[853];
    assign inter_3[854] = inter_2[854];
    assign inter_3[855] = inter_2[855];
    assign inter_3[856] = inter_2[856]^inter_2[860];
    assign inter_3[857] = inter_2[857]^inter_2[861];
    assign inter_3[858] = inter_2[858]^inter_2[862];
    assign inter_3[859] = inter_2[859]^inter_2[863];
    assign inter_3[860] = inter_2[860];
    assign inter_3[861] = inter_2[861];
    assign inter_3[862] = inter_2[862];
    assign inter_3[863] = inter_2[863];
    assign inter_3[864] = inter_2[864]^inter_2[868];
    assign inter_3[865] = inter_2[865]^inter_2[869];
    assign inter_3[866] = inter_2[866]^inter_2[870];
    assign inter_3[867] = inter_2[867]^inter_2[871];
    assign inter_3[868] = inter_2[868];
    assign inter_3[869] = inter_2[869];
    assign inter_3[870] = inter_2[870];
    assign inter_3[871] = inter_2[871];
    assign inter_3[872] = inter_2[872]^inter_2[876];
    assign inter_3[873] = inter_2[873]^inter_2[877];
    assign inter_3[874] = inter_2[874]^inter_2[878];
    assign inter_3[875] = inter_2[875]^inter_2[879];
    assign inter_3[876] = inter_2[876];
    assign inter_3[877] = inter_2[877];
    assign inter_3[878] = inter_2[878];
    assign inter_3[879] = inter_2[879];
    assign inter_3[880] = inter_2[880]^inter_2[884];
    assign inter_3[881] = inter_2[881]^inter_2[885];
    assign inter_3[882] = inter_2[882]^inter_2[886];
    assign inter_3[883] = inter_2[883]^inter_2[887];
    assign inter_3[884] = inter_2[884];
    assign inter_3[885] = inter_2[885];
    assign inter_3[886] = inter_2[886];
    assign inter_3[887] = inter_2[887];
    assign inter_3[888] = inter_2[888]^inter_2[892];
    assign inter_3[889] = inter_2[889]^inter_2[893];
    assign inter_3[890] = inter_2[890]^inter_2[894];
    assign inter_3[891] = inter_2[891]^inter_2[895];
    assign inter_3[892] = inter_2[892];
    assign inter_3[893] = inter_2[893];
    assign inter_3[894] = inter_2[894];
    assign inter_3[895] = inter_2[895];
    assign inter_3[896] = inter_2[896]^inter_2[900];
    assign inter_3[897] = inter_2[897]^inter_2[901];
    assign inter_3[898] = inter_2[898]^inter_2[902];
    assign inter_3[899] = inter_2[899]^inter_2[903];
    assign inter_3[900] = inter_2[900];
    assign inter_3[901] = inter_2[901];
    assign inter_3[902] = inter_2[902];
    assign inter_3[903] = inter_2[903];
    assign inter_3[904] = inter_2[904]^inter_2[908];
    assign inter_3[905] = inter_2[905]^inter_2[909];
    assign inter_3[906] = inter_2[906]^inter_2[910];
    assign inter_3[907] = inter_2[907]^inter_2[911];
    assign inter_3[908] = inter_2[908];
    assign inter_3[909] = inter_2[909];
    assign inter_3[910] = inter_2[910];
    assign inter_3[911] = inter_2[911];
    assign inter_3[912] = inter_2[912]^inter_2[916];
    assign inter_3[913] = inter_2[913]^inter_2[917];
    assign inter_3[914] = inter_2[914]^inter_2[918];
    assign inter_3[915] = inter_2[915]^inter_2[919];
    assign inter_3[916] = inter_2[916];
    assign inter_3[917] = inter_2[917];
    assign inter_3[918] = inter_2[918];
    assign inter_3[919] = inter_2[919];
    assign inter_3[920] = inter_2[920]^inter_2[924];
    assign inter_3[921] = inter_2[921]^inter_2[925];
    assign inter_3[922] = inter_2[922]^inter_2[926];
    assign inter_3[923] = inter_2[923]^inter_2[927];
    assign inter_3[924] = inter_2[924];
    assign inter_3[925] = inter_2[925];
    assign inter_3[926] = inter_2[926];
    assign inter_3[927] = inter_2[927];
    assign inter_3[928] = inter_2[928]^inter_2[932];
    assign inter_3[929] = inter_2[929]^inter_2[933];
    assign inter_3[930] = inter_2[930]^inter_2[934];
    assign inter_3[931] = inter_2[931]^inter_2[935];
    assign inter_3[932] = inter_2[932];
    assign inter_3[933] = inter_2[933];
    assign inter_3[934] = inter_2[934];
    assign inter_3[935] = inter_2[935];
    assign inter_3[936] = inter_2[936]^inter_2[940];
    assign inter_3[937] = inter_2[937]^inter_2[941];
    assign inter_3[938] = inter_2[938]^inter_2[942];
    assign inter_3[939] = inter_2[939]^inter_2[943];
    assign inter_3[940] = inter_2[940];
    assign inter_3[941] = inter_2[941];
    assign inter_3[942] = inter_2[942];
    assign inter_3[943] = inter_2[943];
    assign inter_3[944] = inter_2[944]^inter_2[948];
    assign inter_3[945] = inter_2[945]^inter_2[949];
    assign inter_3[946] = inter_2[946]^inter_2[950];
    assign inter_3[947] = inter_2[947]^inter_2[951];
    assign inter_3[948] = inter_2[948];
    assign inter_3[949] = inter_2[949];
    assign inter_3[950] = inter_2[950];
    assign inter_3[951] = inter_2[951];
    assign inter_3[952] = inter_2[952]^inter_2[956];
    assign inter_3[953] = inter_2[953]^inter_2[957];
    assign inter_3[954] = inter_2[954]^inter_2[958];
    assign inter_3[955] = inter_2[955]^inter_2[959];
    assign inter_3[956] = inter_2[956];
    assign inter_3[957] = inter_2[957];
    assign inter_3[958] = inter_2[958];
    assign inter_3[959] = inter_2[959];
    assign inter_3[960] = inter_2[960]^inter_2[964];
    assign inter_3[961] = inter_2[961]^inter_2[965];
    assign inter_3[962] = inter_2[962]^inter_2[966];
    assign inter_3[963] = inter_2[963]^inter_2[967];
    assign inter_3[964] = inter_2[964];
    assign inter_3[965] = inter_2[965];
    assign inter_3[966] = inter_2[966];
    assign inter_3[967] = inter_2[967];
    assign inter_3[968] = inter_2[968]^inter_2[972];
    assign inter_3[969] = inter_2[969]^inter_2[973];
    assign inter_3[970] = inter_2[970]^inter_2[974];
    assign inter_3[971] = inter_2[971]^inter_2[975];
    assign inter_3[972] = inter_2[972];
    assign inter_3[973] = inter_2[973];
    assign inter_3[974] = inter_2[974];
    assign inter_3[975] = inter_2[975];
    assign inter_3[976] = inter_2[976]^inter_2[980];
    assign inter_3[977] = inter_2[977]^inter_2[981];
    assign inter_3[978] = inter_2[978]^inter_2[982];
    assign inter_3[979] = inter_2[979]^inter_2[983];
    assign inter_3[980] = inter_2[980];
    assign inter_3[981] = inter_2[981];
    assign inter_3[982] = inter_2[982];
    assign inter_3[983] = inter_2[983];
    assign inter_3[984] = inter_2[984]^inter_2[988];
    assign inter_3[985] = inter_2[985]^inter_2[989];
    assign inter_3[986] = inter_2[986]^inter_2[990];
    assign inter_3[987] = inter_2[987]^inter_2[991];
    assign inter_3[988] = inter_2[988];
    assign inter_3[989] = inter_2[989];
    assign inter_3[990] = inter_2[990];
    assign inter_3[991] = inter_2[991];
    assign inter_3[992] = inter_2[992]^inter_2[996];
    assign inter_3[993] = inter_2[993]^inter_2[997];
    assign inter_3[994] = inter_2[994]^inter_2[998];
    assign inter_3[995] = inter_2[995]^inter_2[999];
    assign inter_3[996] = inter_2[996];
    assign inter_3[997] = inter_2[997];
    assign inter_3[998] = inter_2[998];
    assign inter_3[999] = inter_2[999];
    assign inter_3[1000] = inter_2[1000]^inter_2[1004];
    assign inter_3[1001] = inter_2[1001]^inter_2[1005];
    assign inter_3[1002] = inter_2[1002]^inter_2[1006];
    assign inter_3[1003] = inter_2[1003]^inter_2[1007];
    assign inter_3[1004] = inter_2[1004];
    assign inter_3[1005] = inter_2[1005];
    assign inter_3[1006] = inter_2[1006];
    assign inter_3[1007] = inter_2[1007];
    assign inter_3[1008] = inter_2[1008]^inter_2[1012];
    assign inter_3[1009] = inter_2[1009]^inter_2[1013];
    assign inter_3[1010] = inter_2[1010]^inter_2[1014];
    assign inter_3[1011] = inter_2[1011]^inter_2[1015];
    assign inter_3[1012] = inter_2[1012];
    assign inter_3[1013] = inter_2[1013];
    assign inter_3[1014] = inter_2[1014];
    assign inter_3[1015] = inter_2[1015];
    assign inter_3[1016] = inter_2[1016]^inter_2[1020];
    assign inter_3[1017] = inter_2[1017]^inter_2[1021];
    assign inter_3[1018] = inter_2[1018]^inter_2[1022];
    assign inter_3[1019] = inter_2[1019]^inter_2[1023];
    assign inter_3[1020] = inter_2[1020];
    assign inter_3[1021] = inter_2[1021];
    assign inter_3[1022] = inter_2[1022];
    assign inter_3[1023] = inter_2[1023];
    /***************************/
    assign inter_4[0] = inter_3[0]^inter_3[8];
    assign inter_4[1] = inter_3[1]^inter_3[9];
    assign inter_4[2] = inter_3[2]^inter_3[10];
    assign inter_4[3] = inter_3[3]^inter_3[11];
    assign inter_4[4] = inter_3[4]^inter_3[12];
    assign inter_4[5] = inter_3[5]^inter_3[13];
    assign inter_4[6] = inter_3[6]^inter_3[14];
    assign inter_4[7] = inter_3[7]^inter_3[15];
    assign inter_4[8] = inter_3[8];
    assign inter_4[9] = inter_3[9];
    assign inter_4[10] = inter_3[10];
    assign inter_4[11] = inter_3[11];
    assign inter_4[12] = inter_3[12];
    assign inter_4[13] = inter_3[13];
    assign inter_4[14] = inter_3[14];
    assign inter_4[15] = inter_3[15];
    assign inter_4[16] = inter_3[16]^inter_3[24];
    assign inter_4[17] = inter_3[17]^inter_3[25];
    assign inter_4[18] = inter_3[18]^inter_3[26];
    assign inter_4[19] = inter_3[19]^inter_3[27];
    assign inter_4[20] = inter_3[20]^inter_3[28];
    assign inter_4[21] = inter_3[21]^inter_3[29];
    assign inter_4[22] = inter_3[22]^inter_3[30];
    assign inter_4[23] = inter_3[23]^inter_3[31];
    assign inter_4[24] = inter_3[24];
    assign inter_4[25] = inter_3[25];
    assign inter_4[26] = inter_3[26];
    assign inter_4[27] = inter_3[27];
    assign inter_4[28] = inter_3[28];
    assign inter_4[29] = inter_3[29];
    assign inter_4[30] = inter_3[30];
    assign inter_4[31] = inter_3[31];
    assign inter_4[32] = inter_3[32]^inter_3[40];
    assign inter_4[33] = inter_3[33]^inter_3[41];
    assign inter_4[34] = inter_3[34]^inter_3[42];
    assign inter_4[35] = inter_3[35]^inter_3[43];
    assign inter_4[36] = inter_3[36]^inter_3[44];
    assign inter_4[37] = inter_3[37]^inter_3[45];
    assign inter_4[38] = inter_3[38]^inter_3[46];
    assign inter_4[39] = inter_3[39]^inter_3[47];
    assign inter_4[40] = inter_3[40];
    assign inter_4[41] = inter_3[41];
    assign inter_4[42] = inter_3[42];
    assign inter_4[43] = inter_3[43];
    assign inter_4[44] = inter_3[44];
    assign inter_4[45] = inter_3[45];
    assign inter_4[46] = inter_3[46];
    assign inter_4[47] = inter_3[47];
    assign inter_4[48] = inter_3[48]^inter_3[56];
    assign inter_4[49] = inter_3[49]^inter_3[57];
    assign inter_4[50] = inter_3[50]^inter_3[58];
    assign inter_4[51] = inter_3[51]^inter_3[59];
    assign inter_4[52] = inter_3[52]^inter_3[60];
    assign inter_4[53] = inter_3[53]^inter_3[61];
    assign inter_4[54] = inter_3[54]^inter_3[62];
    assign inter_4[55] = inter_3[55]^inter_3[63];
    assign inter_4[56] = inter_3[56];
    assign inter_4[57] = inter_3[57];
    assign inter_4[58] = inter_3[58];
    assign inter_4[59] = inter_3[59];
    assign inter_4[60] = inter_3[60];
    assign inter_4[61] = inter_3[61];
    assign inter_4[62] = inter_3[62];
    assign inter_4[63] = inter_3[63];
    assign inter_4[64] = inter_3[64]^inter_3[72];
    assign inter_4[65] = inter_3[65]^inter_3[73];
    assign inter_4[66] = inter_3[66]^inter_3[74];
    assign inter_4[67] = inter_3[67]^inter_3[75];
    assign inter_4[68] = inter_3[68]^inter_3[76];
    assign inter_4[69] = inter_3[69]^inter_3[77];
    assign inter_4[70] = inter_3[70]^inter_3[78];
    assign inter_4[71] = inter_3[71]^inter_3[79];
    assign inter_4[72] = inter_3[72];
    assign inter_4[73] = inter_3[73];
    assign inter_4[74] = inter_3[74];
    assign inter_4[75] = inter_3[75];
    assign inter_4[76] = inter_3[76];
    assign inter_4[77] = inter_3[77];
    assign inter_4[78] = inter_3[78];
    assign inter_4[79] = inter_3[79];
    assign inter_4[80] = inter_3[80]^inter_3[88];
    assign inter_4[81] = inter_3[81]^inter_3[89];
    assign inter_4[82] = inter_3[82]^inter_3[90];
    assign inter_4[83] = inter_3[83]^inter_3[91];
    assign inter_4[84] = inter_3[84]^inter_3[92];
    assign inter_4[85] = inter_3[85]^inter_3[93];
    assign inter_4[86] = inter_3[86]^inter_3[94];
    assign inter_4[87] = inter_3[87]^inter_3[95];
    assign inter_4[88] = inter_3[88];
    assign inter_4[89] = inter_3[89];
    assign inter_4[90] = inter_3[90];
    assign inter_4[91] = inter_3[91];
    assign inter_4[92] = inter_3[92];
    assign inter_4[93] = inter_3[93];
    assign inter_4[94] = inter_3[94];
    assign inter_4[95] = inter_3[95];
    assign inter_4[96] = inter_3[96]^inter_3[104];
    assign inter_4[97] = inter_3[97]^inter_3[105];
    assign inter_4[98] = inter_3[98]^inter_3[106];
    assign inter_4[99] = inter_3[99]^inter_3[107];
    assign inter_4[100] = inter_3[100]^inter_3[108];
    assign inter_4[101] = inter_3[101]^inter_3[109];
    assign inter_4[102] = inter_3[102]^inter_3[110];
    assign inter_4[103] = inter_3[103]^inter_3[111];
    assign inter_4[104] = inter_3[104];
    assign inter_4[105] = inter_3[105];
    assign inter_4[106] = inter_3[106];
    assign inter_4[107] = inter_3[107];
    assign inter_4[108] = inter_3[108];
    assign inter_4[109] = inter_3[109];
    assign inter_4[110] = inter_3[110];
    assign inter_4[111] = inter_3[111];
    assign inter_4[112] = inter_3[112]^inter_3[120];
    assign inter_4[113] = inter_3[113]^inter_3[121];
    assign inter_4[114] = inter_3[114]^inter_3[122];
    assign inter_4[115] = inter_3[115]^inter_3[123];
    assign inter_4[116] = inter_3[116]^inter_3[124];
    assign inter_4[117] = inter_3[117]^inter_3[125];
    assign inter_4[118] = inter_3[118]^inter_3[126];
    assign inter_4[119] = inter_3[119]^inter_3[127];
    assign inter_4[120] = inter_3[120];
    assign inter_4[121] = inter_3[121];
    assign inter_4[122] = inter_3[122];
    assign inter_4[123] = inter_3[123];
    assign inter_4[124] = inter_3[124];
    assign inter_4[125] = inter_3[125];
    assign inter_4[126] = inter_3[126];
    assign inter_4[127] = inter_3[127];
    assign inter_4[128] = inter_3[128]^inter_3[136];
    assign inter_4[129] = inter_3[129]^inter_3[137];
    assign inter_4[130] = inter_3[130]^inter_3[138];
    assign inter_4[131] = inter_3[131]^inter_3[139];
    assign inter_4[132] = inter_3[132]^inter_3[140];
    assign inter_4[133] = inter_3[133]^inter_3[141];
    assign inter_4[134] = inter_3[134]^inter_3[142];
    assign inter_4[135] = inter_3[135]^inter_3[143];
    assign inter_4[136] = inter_3[136];
    assign inter_4[137] = inter_3[137];
    assign inter_4[138] = inter_3[138];
    assign inter_4[139] = inter_3[139];
    assign inter_4[140] = inter_3[140];
    assign inter_4[141] = inter_3[141];
    assign inter_4[142] = inter_3[142];
    assign inter_4[143] = inter_3[143];
    assign inter_4[144] = inter_3[144]^inter_3[152];
    assign inter_4[145] = inter_3[145]^inter_3[153];
    assign inter_4[146] = inter_3[146]^inter_3[154];
    assign inter_4[147] = inter_3[147]^inter_3[155];
    assign inter_4[148] = inter_3[148]^inter_3[156];
    assign inter_4[149] = inter_3[149]^inter_3[157];
    assign inter_4[150] = inter_3[150]^inter_3[158];
    assign inter_4[151] = inter_3[151]^inter_3[159];
    assign inter_4[152] = inter_3[152];
    assign inter_4[153] = inter_3[153];
    assign inter_4[154] = inter_3[154];
    assign inter_4[155] = inter_3[155];
    assign inter_4[156] = inter_3[156];
    assign inter_4[157] = inter_3[157];
    assign inter_4[158] = inter_3[158];
    assign inter_4[159] = inter_3[159];
    assign inter_4[160] = inter_3[160]^inter_3[168];
    assign inter_4[161] = inter_3[161]^inter_3[169];
    assign inter_4[162] = inter_3[162]^inter_3[170];
    assign inter_4[163] = inter_3[163]^inter_3[171];
    assign inter_4[164] = inter_3[164]^inter_3[172];
    assign inter_4[165] = inter_3[165]^inter_3[173];
    assign inter_4[166] = inter_3[166]^inter_3[174];
    assign inter_4[167] = inter_3[167]^inter_3[175];
    assign inter_4[168] = inter_3[168];
    assign inter_4[169] = inter_3[169];
    assign inter_4[170] = inter_3[170];
    assign inter_4[171] = inter_3[171];
    assign inter_4[172] = inter_3[172];
    assign inter_4[173] = inter_3[173];
    assign inter_4[174] = inter_3[174];
    assign inter_4[175] = inter_3[175];
    assign inter_4[176] = inter_3[176]^inter_3[184];
    assign inter_4[177] = inter_3[177]^inter_3[185];
    assign inter_4[178] = inter_3[178]^inter_3[186];
    assign inter_4[179] = inter_3[179]^inter_3[187];
    assign inter_4[180] = inter_3[180]^inter_3[188];
    assign inter_4[181] = inter_3[181]^inter_3[189];
    assign inter_4[182] = inter_3[182]^inter_3[190];
    assign inter_4[183] = inter_3[183]^inter_3[191];
    assign inter_4[184] = inter_3[184];
    assign inter_4[185] = inter_3[185];
    assign inter_4[186] = inter_3[186];
    assign inter_4[187] = inter_3[187];
    assign inter_4[188] = inter_3[188];
    assign inter_4[189] = inter_3[189];
    assign inter_4[190] = inter_3[190];
    assign inter_4[191] = inter_3[191];
    assign inter_4[192] = inter_3[192]^inter_3[200];
    assign inter_4[193] = inter_3[193]^inter_3[201];
    assign inter_4[194] = inter_3[194]^inter_3[202];
    assign inter_4[195] = inter_3[195]^inter_3[203];
    assign inter_4[196] = inter_3[196]^inter_3[204];
    assign inter_4[197] = inter_3[197]^inter_3[205];
    assign inter_4[198] = inter_3[198]^inter_3[206];
    assign inter_4[199] = inter_3[199]^inter_3[207];
    assign inter_4[200] = inter_3[200];
    assign inter_4[201] = inter_3[201];
    assign inter_4[202] = inter_3[202];
    assign inter_4[203] = inter_3[203];
    assign inter_4[204] = inter_3[204];
    assign inter_4[205] = inter_3[205];
    assign inter_4[206] = inter_3[206];
    assign inter_4[207] = inter_3[207];
    assign inter_4[208] = inter_3[208]^inter_3[216];
    assign inter_4[209] = inter_3[209]^inter_3[217];
    assign inter_4[210] = inter_3[210]^inter_3[218];
    assign inter_4[211] = inter_3[211]^inter_3[219];
    assign inter_4[212] = inter_3[212]^inter_3[220];
    assign inter_4[213] = inter_3[213]^inter_3[221];
    assign inter_4[214] = inter_3[214]^inter_3[222];
    assign inter_4[215] = inter_3[215]^inter_3[223];
    assign inter_4[216] = inter_3[216];
    assign inter_4[217] = inter_3[217];
    assign inter_4[218] = inter_3[218];
    assign inter_4[219] = inter_3[219];
    assign inter_4[220] = inter_3[220];
    assign inter_4[221] = inter_3[221];
    assign inter_4[222] = inter_3[222];
    assign inter_4[223] = inter_3[223];
    assign inter_4[224] = inter_3[224]^inter_3[232];
    assign inter_4[225] = inter_3[225]^inter_3[233];
    assign inter_4[226] = inter_3[226]^inter_3[234];
    assign inter_4[227] = inter_3[227]^inter_3[235];
    assign inter_4[228] = inter_3[228]^inter_3[236];
    assign inter_4[229] = inter_3[229]^inter_3[237];
    assign inter_4[230] = inter_3[230]^inter_3[238];
    assign inter_4[231] = inter_3[231]^inter_3[239];
    assign inter_4[232] = inter_3[232];
    assign inter_4[233] = inter_3[233];
    assign inter_4[234] = inter_3[234];
    assign inter_4[235] = inter_3[235];
    assign inter_4[236] = inter_3[236];
    assign inter_4[237] = inter_3[237];
    assign inter_4[238] = inter_3[238];
    assign inter_4[239] = inter_3[239];
    assign inter_4[240] = inter_3[240]^inter_3[248];
    assign inter_4[241] = inter_3[241]^inter_3[249];
    assign inter_4[242] = inter_3[242]^inter_3[250];
    assign inter_4[243] = inter_3[243]^inter_3[251];
    assign inter_4[244] = inter_3[244]^inter_3[252];
    assign inter_4[245] = inter_3[245]^inter_3[253];
    assign inter_4[246] = inter_3[246]^inter_3[254];
    assign inter_4[247] = inter_3[247]^inter_3[255];
    assign inter_4[248] = inter_3[248];
    assign inter_4[249] = inter_3[249];
    assign inter_4[250] = inter_3[250];
    assign inter_4[251] = inter_3[251];
    assign inter_4[252] = inter_3[252];
    assign inter_4[253] = inter_3[253];
    assign inter_4[254] = inter_3[254];
    assign inter_4[255] = inter_3[255];
    assign inter_4[256] = inter_3[256]^inter_3[264];
    assign inter_4[257] = inter_3[257]^inter_3[265];
    assign inter_4[258] = inter_3[258]^inter_3[266];
    assign inter_4[259] = inter_3[259]^inter_3[267];
    assign inter_4[260] = inter_3[260]^inter_3[268];
    assign inter_4[261] = inter_3[261]^inter_3[269];
    assign inter_4[262] = inter_3[262]^inter_3[270];
    assign inter_4[263] = inter_3[263]^inter_3[271];
    assign inter_4[264] = inter_3[264];
    assign inter_4[265] = inter_3[265];
    assign inter_4[266] = inter_3[266];
    assign inter_4[267] = inter_3[267];
    assign inter_4[268] = inter_3[268];
    assign inter_4[269] = inter_3[269];
    assign inter_4[270] = inter_3[270];
    assign inter_4[271] = inter_3[271];
    assign inter_4[272] = inter_3[272]^inter_3[280];
    assign inter_4[273] = inter_3[273]^inter_3[281];
    assign inter_4[274] = inter_3[274]^inter_3[282];
    assign inter_4[275] = inter_3[275]^inter_3[283];
    assign inter_4[276] = inter_3[276]^inter_3[284];
    assign inter_4[277] = inter_3[277]^inter_3[285];
    assign inter_4[278] = inter_3[278]^inter_3[286];
    assign inter_4[279] = inter_3[279]^inter_3[287];
    assign inter_4[280] = inter_3[280];
    assign inter_4[281] = inter_3[281];
    assign inter_4[282] = inter_3[282];
    assign inter_4[283] = inter_3[283];
    assign inter_4[284] = inter_3[284];
    assign inter_4[285] = inter_3[285];
    assign inter_4[286] = inter_3[286];
    assign inter_4[287] = inter_3[287];
    assign inter_4[288] = inter_3[288]^inter_3[296];
    assign inter_4[289] = inter_3[289]^inter_3[297];
    assign inter_4[290] = inter_3[290]^inter_3[298];
    assign inter_4[291] = inter_3[291]^inter_3[299];
    assign inter_4[292] = inter_3[292]^inter_3[300];
    assign inter_4[293] = inter_3[293]^inter_3[301];
    assign inter_4[294] = inter_3[294]^inter_3[302];
    assign inter_4[295] = inter_3[295]^inter_3[303];
    assign inter_4[296] = inter_3[296];
    assign inter_4[297] = inter_3[297];
    assign inter_4[298] = inter_3[298];
    assign inter_4[299] = inter_3[299];
    assign inter_4[300] = inter_3[300];
    assign inter_4[301] = inter_3[301];
    assign inter_4[302] = inter_3[302];
    assign inter_4[303] = inter_3[303];
    assign inter_4[304] = inter_3[304]^inter_3[312];
    assign inter_4[305] = inter_3[305]^inter_3[313];
    assign inter_4[306] = inter_3[306]^inter_3[314];
    assign inter_4[307] = inter_3[307]^inter_3[315];
    assign inter_4[308] = inter_3[308]^inter_3[316];
    assign inter_4[309] = inter_3[309]^inter_3[317];
    assign inter_4[310] = inter_3[310]^inter_3[318];
    assign inter_4[311] = inter_3[311]^inter_3[319];
    assign inter_4[312] = inter_3[312];
    assign inter_4[313] = inter_3[313];
    assign inter_4[314] = inter_3[314];
    assign inter_4[315] = inter_3[315];
    assign inter_4[316] = inter_3[316];
    assign inter_4[317] = inter_3[317];
    assign inter_4[318] = inter_3[318];
    assign inter_4[319] = inter_3[319];
    assign inter_4[320] = inter_3[320]^inter_3[328];
    assign inter_4[321] = inter_3[321]^inter_3[329];
    assign inter_4[322] = inter_3[322]^inter_3[330];
    assign inter_4[323] = inter_3[323]^inter_3[331];
    assign inter_4[324] = inter_3[324]^inter_3[332];
    assign inter_4[325] = inter_3[325]^inter_3[333];
    assign inter_4[326] = inter_3[326]^inter_3[334];
    assign inter_4[327] = inter_3[327]^inter_3[335];
    assign inter_4[328] = inter_3[328];
    assign inter_4[329] = inter_3[329];
    assign inter_4[330] = inter_3[330];
    assign inter_4[331] = inter_3[331];
    assign inter_4[332] = inter_3[332];
    assign inter_4[333] = inter_3[333];
    assign inter_4[334] = inter_3[334];
    assign inter_4[335] = inter_3[335];
    assign inter_4[336] = inter_3[336]^inter_3[344];
    assign inter_4[337] = inter_3[337]^inter_3[345];
    assign inter_4[338] = inter_3[338]^inter_3[346];
    assign inter_4[339] = inter_3[339]^inter_3[347];
    assign inter_4[340] = inter_3[340]^inter_3[348];
    assign inter_4[341] = inter_3[341]^inter_3[349];
    assign inter_4[342] = inter_3[342]^inter_3[350];
    assign inter_4[343] = inter_3[343]^inter_3[351];
    assign inter_4[344] = inter_3[344];
    assign inter_4[345] = inter_3[345];
    assign inter_4[346] = inter_3[346];
    assign inter_4[347] = inter_3[347];
    assign inter_4[348] = inter_3[348];
    assign inter_4[349] = inter_3[349];
    assign inter_4[350] = inter_3[350];
    assign inter_4[351] = inter_3[351];
    assign inter_4[352] = inter_3[352]^inter_3[360];
    assign inter_4[353] = inter_3[353]^inter_3[361];
    assign inter_4[354] = inter_3[354]^inter_3[362];
    assign inter_4[355] = inter_3[355]^inter_3[363];
    assign inter_4[356] = inter_3[356]^inter_3[364];
    assign inter_4[357] = inter_3[357]^inter_3[365];
    assign inter_4[358] = inter_3[358]^inter_3[366];
    assign inter_4[359] = inter_3[359]^inter_3[367];
    assign inter_4[360] = inter_3[360];
    assign inter_4[361] = inter_3[361];
    assign inter_4[362] = inter_3[362];
    assign inter_4[363] = inter_3[363];
    assign inter_4[364] = inter_3[364];
    assign inter_4[365] = inter_3[365];
    assign inter_4[366] = inter_3[366];
    assign inter_4[367] = inter_3[367];
    assign inter_4[368] = inter_3[368]^inter_3[376];
    assign inter_4[369] = inter_3[369]^inter_3[377];
    assign inter_4[370] = inter_3[370]^inter_3[378];
    assign inter_4[371] = inter_3[371]^inter_3[379];
    assign inter_4[372] = inter_3[372]^inter_3[380];
    assign inter_4[373] = inter_3[373]^inter_3[381];
    assign inter_4[374] = inter_3[374]^inter_3[382];
    assign inter_4[375] = inter_3[375]^inter_3[383];
    assign inter_4[376] = inter_3[376];
    assign inter_4[377] = inter_3[377];
    assign inter_4[378] = inter_3[378];
    assign inter_4[379] = inter_3[379];
    assign inter_4[380] = inter_3[380];
    assign inter_4[381] = inter_3[381];
    assign inter_4[382] = inter_3[382];
    assign inter_4[383] = inter_3[383];
    assign inter_4[384] = inter_3[384]^inter_3[392];
    assign inter_4[385] = inter_3[385]^inter_3[393];
    assign inter_4[386] = inter_3[386]^inter_3[394];
    assign inter_4[387] = inter_3[387]^inter_3[395];
    assign inter_4[388] = inter_3[388]^inter_3[396];
    assign inter_4[389] = inter_3[389]^inter_3[397];
    assign inter_4[390] = inter_3[390]^inter_3[398];
    assign inter_4[391] = inter_3[391]^inter_3[399];
    assign inter_4[392] = inter_3[392];
    assign inter_4[393] = inter_3[393];
    assign inter_4[394] = inter_3[394];
    assign inter_4[395] = inter_3[395];
    assign inter_4[396] = inter_3[396];
    assign inter_4[397] = inter_3[397];
    assign inter_4[398] = inter_3[398];
    assign inter_4[399] = inter_3[399];
    assign inter_4[400] = inter_3[400]^inter_3[408];
    assign inter_4[401] = inter_3[401]^inter_3[409];
    assign inter_4[402] = inter_3[402]^inter_3[410];
    assign inter_4[403] = inter_3[403]^inter_3[411];
    assign inter_4[404] = inter_3[404]^inter_3[412];
    assign inter_4[405] = inter_3[405]^inter_3[413];
    assign inter_4[406] = inter_3[406]^inter_3[414];
    assign inter_4[407] = inter_3[407]^inter_3[415];
    assign inter_4[408] = inter_3[408];
    assign inter_4[409] = inter_3[409];
    assign inter_4[410] = inter_3[410];
    assign inter_4[411] = inter_3[411];
    assign inter_4[412] = inter_3[412];
    assign inter_4[413] = inter_3[413];
    assign inter_4[414] = inter_3[414];
    assign inter_4[415] = inter_3[415];
    assign inter_4[416] = inter_3[416]^inter_3[424];
    assign inter_4[417] = inter_3[417]^inter_3[425];
    assign inter_4[418] = inter_3[418]^inter_3[426];
    assign inter_4[419] = inter_3[419]^inter_3[427];
    assign inter_4[420] = inter_3[420]^inter_3[428];
    assign inter_4[421] = inter_3[421]^inter_3[429];
    assign inter_4[422] = inter_3[422]^inter_3[430];
    assign inter_4[423] = inter_3[423]^inter_3[431];
    assign inter_4[424] = inter_3[424];
    assign inter_4[425] = inter_3[425];
    assign inter_4[426] = inter_3[426];
    assign inter_4[427] = inter_3[427];
    assign inter_4[428] = inter_3[428];
    assign inter_4[429] = inter_3[429];
    assign inter_4[430] = inter_3[430];
    assign inter_4[431] = inter_3[431];
    assign inter_4[432] = inter_3[432]^inter_3[440];
    assign inter_4[433] = inter_3[433]^inter_3[441];
    assign inter_4[434] = inter_3[434]^inter_3[442];
    assign inter_4[435] = inter_3[435]^inter_3[443];
    assign inter_4[436] = inter_3[436]^inter_3[444];
    assign inter_4[437] = inter_3[437]^inter_3[445];
    assign inter_4[438] = inter_3[438]^inter_3[446];
    assign inter_4[439] = inter_3[439]^inter_3[447];
    assign inter_4[440] = inter_3[440];
    assign inter_4[441] = inter_3[441];
    assign inter_4[442] = inter_3[442];
    assign inter_4[443] = inter_3[443];
    assign inter_4[444] = inter_3[444];
    assign inter_4[445] = inter_3[445];
    assign inter_4[446] = inter_3[446];
    assign inter_4[447] = inter_3[447];
    assign inter_4[448] = inter_3[448]^inter_3[456];
    assign inter_4[449] = inter_3[449]^inter_3[457];
    assign inter_4[450] = inter_3[450]^inter_3[458];
    assign inter_4[451] = inter_3[451]^inter_3[459];
    assign inter_4[452] = inter_3[452]^inter_3[460];
    assign inter_4[453] = inter_3[453]^inter_3[461];
    assign inter_4[454] = inter_3[454]^inter_3[462];
    assign inter_4[455] = inter_3[455]^inter_3[463];
    assign inter_4[456] = inter_3[456];
    assign inter_4[457] = inter_3[457];
    assign inter_4[458] = inter_3[458];
    assign inter_4[459] = inter_3[459];
    assign inter_4[460] = inter_3[460];
    assign inter_4[461] = inter_3[461];
    assign inter_4[462] = inter_3[462];
    assign inter_4[463] = inter_3[463];
    assign inter_4[464] = inter_3[464]^inter_3[472];
    assign inter_4[465] = inter_3[465]^inter_3[473];
    assign inter_4[466] = inter_3[466]^inter_3[474];
    assign inter_4[467] = inter_3[467]^inter_3[475];
    assign inter_4[468] = inter_3[468]^inter_3[476];
    assign inter_4[469] = inter_3[469]^inter_3[477];
    assign inter_4[470] = inter_3[470]^inter_3[478];
    assign inter_4[471] = inter_3[471]^inter_3[479];
    assign inter_4[472] = inter_3[472];
    assign inter_4[473] = inter_3[473];
    assign inter_4[474] = inter_3[474];
    assign inter_4[475] = inter_3[475];
    assign inter_4[476] = inter_3[476];
    assign inter_4[477] = inter_3[477];
    assign inter_4[478] = inter_3[478];
    assign inter_4[479] = inter_3[479];
    assign inter_4[480] = inter_3[480]^inter_3[488];
    assign inter_4[481] = inter_3[481]^inter_3[489];
    assign inter_4[482] = inter_3[482]^inter_3[490];
    assign inter_4[483] = inter_3[483]^inter_3[491];
    assign inter_4[484] = inter_3[484]^inter_3[492];
    assign inter_4[485] = inter_3[485]^inter_3[493];
    assign inter_4[486] = inter_3[486]^inter_3[494];
    assign inter_4[487] = inter_3[487]^inter_3[495];
    assign inter_4[488] = inter_3[488];
    assign inter_4[489] = inter_3[489];
    assign inter_4[490] = inter_3[490];
    assign inter_4[491] = inter_3[491];
    assign inter_4[492] = inter_3[492];
    assign inter_4[493] = inter_3[493];
    assign inter_4[494] = inter_3[494];
    assign inter_4[495] = inter_3[495];
    assign inter_4[496] = inter_3[496]^inter_3[504];
    assign inter_4[497] = inter_3[497]^inter_3[505];
    assign inter_4[498] = inter_3[498]^inter_3[506];
    assign inter_4[499] = inter_3[499]^inter_3[507];
    assign inter_4[500] = inter_3[500]^inter_3[508];
    assign inter_4[501] = inter_3[501]^inter_3[509];
    assign inter_4[502] = inter_3[502]^inter_3[510];
    assign inter_4[503] = inter_3[503]^inter_3[511];
    assign inter_4[504] = inter_3[504];
    assign inter_4[505] = inter_3[505];
    assign inter_4[506] = inter_3[506];
    assign inter_4[507] = inter_3[507];
    assign inter_4[508] = inter_3[508];
    assign inter_4[509] = inter_3[509];
    assign inter_4[510] = inter_3[510];
    assign inter_4[511] = inter_3[511];
    assign inter_4[512] = inter_3[512]^inter_3[520];
    assign inter_4[513] = inter_3[513]^inter_3[521];
    assign inter_4[514] = inter_3[514]^inter_3[522];
    assign inter_4[515] = inter_3[515]^inter_3[523];
    assign inter_4[516] = inter_3[516]^inter_3[524];
    assign inter_4[517] = inter_3[517]^inter_3[525];
    assign inter_4[518] = inter_3[518]^inter_3[526];
    assign inter_4[519] = inter_3[519]^inter_3[527];
    assign inter_4[520] = inter_3[520];
    assign inter_4[521] = inter_3[521];
    assign inter_4[522] = inter_3[522];
    assign inter_4[523] = inter_3[523];
    assign inter_4[524] = inter_3[524];
    assign inter_4[525] = inter_3[525];
    assign inter_4[526] = inter_3[526];
    assign inter_4[527] = inter_3[527];
    assign inter_4[528] = inter_3[528]^inter_3[536];
    assign inter_4[529] = inter_3[529]^inter_3[537];
    assign inter_4[530] = inter_3[530]^inter_3[538];
    assign inter_4[531] = inter_3[531]^inter_3[539];
    assign inter_4[532] = inter_3[532]^inter_3[540];
    assign inter_4[533] = inter_3[533]^inter_3[541];
    assign inter_4[534] = inter_3[534]^inter_3[542];
    assign inter_4[535] = inter_3[535]^inter_3[543];
    assign inter_4[536] = inter_3[536];
    assign inter_4[537] = inter_3[537];
    assign inter_4[538] = inter_3[538];
    assign inter_4[539] = inter_3[539];
    assign inter_4[540] = inter_3[540];
    assign inter_4[541] = inter_3[541];
    assign inter_4[542] = inter_3[542];
    assign inter_4[543] = inter_3[543];
    assign inter_4[544] = inter_3[544]^inter_3[552];
    assign inter_4[545] = inter_3[545]^inter_3[553];
    assign inter_4[546] = inter_3[546]^inter_3[554];
    assign inter_4[547] = inter_3[547]^inter_3[555];
    assign inter_4[548] = inter_3[548]^inter_3[556];
    assign inter_4[549] = inter_3[549]^inter_3[557];
    assign inter_4[550] = inter_3[550]^inter_3[558];
    assign inter_4[551] = inter_3[551]^inter_3[559];
    assign inter_4[552] = inter_3[552];
    assign inter_4[553] = inter_3[553];
    assign inter_4[554] = inter_3[554];
    assign inter_4[555] = inter_3[555];
    assign inter_4[556] = inter_3[556];
    assign inter_4[557] = inter_3[557];
    assign inter_4[558] = inter_3[558];
    assign inter_4[559] = inter_3[559];
    assign inter_4[560] = inter_3[560]^inter_3[568];
    assign inter_4[561] = inter_3[561]^inter_3[569];
    assign inter_4[562] = inter_3[562]^inter_3[570];
    assign inter_4[563] = inter_3[563]^inter_3[571];
    assign inter_4[564] = inter_3[564]^inter_3[572];
    assign inter_4[565] = inter_3[565]^inter_3[573];
    assign inter_4[566] = inter_3[566]^inter_3[574];
    assign inter_4[567] = inter_3[567]^inter_3[575];
    assign inter_4[568] = inter_3[568];
    assign inter_4[569] = inter_3[569];
    assign inter_4[570] = inter_3[570];
    assign inter_4[571] = inter_3[571];
    assign inter_4[572] = inter_3[572];
    assign inter_4[573] = inter_3[573];
    assign inter_4[574] = inter_3[574];
    assign inter_4[575] = inter_3[575];
    assign inter_4[576] = inter_3[576]^inter_3[584];
    assign inter_4[577] = inter_3[577]^inter_3[585];
    assign inter_4[578] = inter_3[578]^inter_3[586];
    assign inter_4[579] = inter_3[579]^inter_3[587];
    assign inter_4[580] = inter_3[580]^inter_3[588];
    assign inter_4[581] = inter_3[581]^inter_3[589];
    assign inter_4[582] = inter_3[582]^inter_3[590];
    assign inter_4[583] = inter_3[583]^inter_3[591];
    assign inter_4[584] = inter_3[584];
    assign inter_4[585] = inter_3[585];
    assign inter_4[586] = inter_3[586];
    assign inter_4[587] = inter_3[587];
    assign inter_4[588] = inter_3[588];
    assign inter_4[589] = inter_3[589];
    assign inter_4[590] = inter_3[590];
    assign inter_4[591] = inter_3[591];
    assign inter_4[592] = inter_3[592]^inter_3[600];
    assign inter_4[593] = inter_3[593]^inter_3[601];
    assign inter_4[594] = inter_3[594]^inter_3[602];
    assign inter_4[595] = inter_3[595]^inter_3[603];
    assign inter_4[596] = inter_3[596]^inter_3[604];
    assign inter_4[597] = inter_3[597]^inter_3[605];
    assign inter_4[598] = inter_3[598]^inter_3[606];
    assign inter_4[599] = inter_3[599]^inter_3[607];
    assign inter_4[600] = inter_3[600];
    assign inter_4[601] = inter_3[601];
    assign inter_4[602] = inter_3[602];
    assign inter_4[603] = inter_3[603];
    assign inter_4[604] = inter_3[604];
    assign inter_4[605] = inter_3[605];
    assign inter_4[606] = inter_3[606];
    assign inter_4[607] = inter_3[607];
    assign inter_4[608] = inter_3[608]^inter_3[616];
    assign inter_4[609] = inter_3[609]^inter_3[617];
    assign inter_4[610] = inter_3[610]^inter_3[618];
    assign inter_4[611] = inter_3[611]^inter_3[619];
    assign inter_4[612] = inter_3[612]^inter_3[620];
    assign inter_4[613] = inter_3[613]^inter_3[621];
    assign inter_4[614] = inter_3[614]^inter_3[622];
    assign inter_4[615] = inter_3[615]^inter_3[623];
    assign inter_4[616] = inter_3[616];
    assign inter_4[617] = inter_3[617];
    assign inter_4[618] = inter_3[618];
    assign inter_4[619] = inter_3[619];
    assign inter_4[620] = inter_3[620];
    assign inter_4[621] = inter_3[621];
    assign inter_4[622] = inter_3[622];
    assign inter_4[623] = inter_3[623];
    assign inter_4[624] = inter_3[624]^inter_3[632];
    assign inter_4[625] = inter_3[625]^inter_3[633];
    assign inter_4[626] = inter_3[626]^inter_3[634];
    assign inter_4[627] = inter_3[627]^inter_3[635];
    assign inter_4[628] = inter_3[628]^inter_3[636];
    assign inter_4[629] = inter_3[629]^inter_3[637];
    assign inter_4[630] = inter_3[630]^inter_3[638];
    assign inter_4[631] = inter_3[631]^inter_3[639];
    assign inter_4[632] = inter_3[632];
    assign inter_4[633] = inter_3[633];
    assign inter_4[634] = inter_3[634];
    assign inter_4[635] = inter_3[635];
    assign inter_4[636] = inter_3[636];
    assign inter_4[637] = inter_3[637];
    assign inter_4[638] = inter_3[638];
    assign inter_4[639] = inter_3[639];
    assign inter_4[640] = inter_3[640]^inter_3[648];
    assign inter_4[641] = inter_3[641]^inter_3[649];
    assign inter_4[642] = inter_3[642]^inter_3[650];
    assign inter_4[643] = inter_3[643]^inter_3[651];
    assign inter_4[644] = inter_3[644]^inter_3[652];
    assign inter_4[645] = inter_3[645]^inter_3[653];
    assign inter_4[646] = inter_3[646]^inter_3[654];
    assign inter_4[647] = inter_3[647]^inter_3[655];
    assign inter_4[648] = inter_3[648];
    assign inter_4[649] = inter_3[649];
    assign inter_4[650] = inter_3[650];
    assign inter_4[651] = inter_3[651];
    assign inter_4[652] = inter_3[652];
    assign inter_4[653] = inter_3[653];
    assign inter_4[654] = inter_3[654];
    assign inter_4[655] = inter_3[655];
    assign inter_4[656] = inter_3[656]^inter_3[664];
    assign inter_4[657] = inter_3[657]^inter_3[665];
    assign inter_4[658] = inter_3[658]^inter_3[666];
    assign inter_4[659] = inter_3[659]^inter_3[667];
    assign inter_4[660] = inter_3[660]^inter_3[668];
    assign inter_4[661] = inter_3[661]^inter_3[669];
    assign inter_4[662] = inter_3[662]^inter_3[670];
    assign inter_4[663] = inter_3[663]^inter_3[671];
    assign inter_4[664] = inter_3[664];
    assign inter_4[665] = inter_3[665];
    assign inter_4[666] = inter_3[666];
    assign inter_4[667] = inter_3[667];
    assign inter_4[668] = inter_3[668];
    assign inter_4[669] = inter_3[669];
    assign inter_4[670] = inter_3[670];
    assign inter_4[671] = inter_3[671];
    assign inter_4[672] = inter_3[672]^inter_3[680];
    assign inter_4[673] = inter_3[673]^inter_3[681];
    assign inter_4[674] = inter_3[674]^inter_3[682];
    assign inter_4[675] = inter_3[675]^inter_3[683];
    assign inter_4[676] = inter_3[676]^inter_3[684];
    assign inter_4[677] = inter_3[677]^inter_3[685];
    assign inter_4[678] = inter_3[678]^inter_3[686];
    assign inter_4[679] = inter_3[679]^inter_3[687];
    assign inter_4[680] = inter_3[680];
    assign inter_4[681] = inter_3[681];
    assign inter_4[682] = inter_3[682];
    assign inter_4[683] = inter_3[683];
    assign inter_4[684] = inter_3[684];
    assign inter_4[685] = inter_3[685];
    assign inter_4[686] = inter_3[686];
    assign inter_4[687] = inter_3[687];
    assign inter_4[688] = inter_3[688]^inter_3[696];
    assign inter_4[689] = inter_3[689]^inter_3[697];
    assign inter_4[690] = inter_3[690]^inter_3[698];
    assign inter_4[691] = inter_3[691]^inter_3[699];
    assign inter_4[692] = inter_3[692]^inter_3[700];
    assign inter_4[693] = inter_3[693]^inter_3[701];
    assign inter_4[694] = inter_3[694]^inter_3[702];
    assign inter_4[695] = inter_3[695]^inter_3[703];
    assign inter_4[696] = inter_3[696];
    assign inter_4[697] = inter_3[697];
    assign inter_4[698] = inter_3[698];
    assign inter_4[699] = inter_3[699];
    assign inter_4[700] = inter_3[700];
    assign inter_4[701] = inter_3[701];
    assign inter_4[702] = inter_3[702];
    assign inter_4[703] = inter_3[703];
    assign inter_4[704] = inter_3[704]^inter_3[712];
    assign inter_4[705] = inter_3[705]^inter_3[713];
    assign inter_4[706] = inter_3[706]^inter_3[714];
    assign inter_4[707] = inter_3[707]^inter_3[715];
    assign inter_4[708] = inter_3[708]^inter_3[716];
    assign inter_4[709] = inter_3[709]^inter_3[717];
    assign inter_4[710] = inter_3[710]^inter_3[718];
    assign inter_4[711] = inter_3[711]^inter_3[719];
    assign inter_4[712] = inter_3[712];
    assign inter_4[713] = inter_3[713];
    assign inter_4[714] = inter_3[714];
    assign inter_4[715] = inter_3[715];
    assign inter_4[716] = inter_3[716];
    assign inter_4[717] = inter_3[717];
    assign inter_4[718] = inter_3[718];
    assign inter_4[719] = inter_3[719];
    assign inter_4[720] = inter_3[720]^inter_3[728];
    assign inter_4[721] = inter_3[721]^inter_3[729];
    assign inter_4[722] = inter_3[722]^inter_3[730];
    assign inter_4[723] = inter_3[723]^inter_3[731];
    assign inter_4[724] = inter_3[724]^inter_3[732];
    assign inter_4[725] = inter_3[725]^inter_3[733];
    assign inter_4[726] = inter_3[726]^inter_3[734];
    assign inter_4[727] = inter_3[727]^inter_3[735];
    assign inter_4[728] = inter_3[728];
    assign inter_4[729] = inter_3[729];
    assign inter_4[730] = inter_3[730];
    assign inter_4[731] = inter_3[731];
    assign inter_4[732] = inter_3[732];
    assign inter_4[733] = inter_3[733];
    assign inter_4[734] = inter_3[734];
    assign inter_4[735] = inter_3[735];
    assign inter_4[736] = inter_3[736]^inter_3[744];
    assign inter_4[737] = inter_3[737]^inter_3[745];
    assign inter_4[738] = inter_3[738]^inter_3[746];
    assign inter_4[739] = inter_3[739]^inter_3[747];
    assign inter_4[740] = inter_3[740]^inter_3[748];
    assign inter_4[741] = inter_3[741]^inter_3[749];
    assign inter_4[742] = inter_3[742]^inter_3[750];
    assign inter_4[743] = inter_3[743]^inter_3[751];
    assign inter_4[744] = inter_3[744];
    assign inter_4[745] = inter_3[745];
    assign inter_4[746] = inter_3[746];
    assign inter_4[747] = inter_3[747];
    assign inter_4[748] = inter_3[748];
    assign inter_4[749] = inter_3[749];
    assign inter_4[750] = inter_3[750];
    assign inter_4[751] = inter_3[751];
    assign inter_4[752] = inter_3[752]^inter_3[760];
    assign inter_4[753] = inter_3[753]^inter_3[761];
    assign inter_4[754] = inter_3[754]^inter_3[762];
    assign inter_4[755] = inter_3[755]^inter_3[763];
    assign inter_4[756] = inter_3[756]^inter_3[764];
    assign inter_4[757] = inter_3[757]^inter_3[765];
    assign inter_4[758] = inter_3[758]^inter_3[766];
    assign inter_4[759] = inter_3[759]^inter_3[767];
    assign inter_4[760] = inter_3[760];
    assign inter_4[761] = inter_3[761];
    assign inter_4[762] = inter_3[762];
    assign inter_4[763] = inter_3[763];
    assign inter_4[764] = inter_3[764];
    assign inter_4[765] = inter_3[765];
    assign inter_4[766] = inter_3[766];
    assign inter_4[767] = inter_3[767];
    assign inter_4[768] = inter_3[768]^inter_3[776];
    assign inter_4[769] = inter_3[769]^inter_3[777];
    assign inter_4[770] = inter_3[770]^inter_3[778];
    assign inter_4[771] = inter_3[771]^inter_3[779];
    assign inter_4[772] = inter_3[772]^inter_3[780];
    assign inter_4[773] = inter_3[773]^inter_3[781];
    assign inter_4[774] = inter_3[774]^inter_3[782];
    assign inter_4[775] = inter_3[775]^inter_3[783];
    assign inter_4[776] = inter_3[776];
    assign inter_4[777] = inter_3[777];
    assign inter_4[778] = inter_3[778];
    assign inter_4[779] = inter_3[779];
    assign inter_4[780] = inter_3[780];
    assign inter_4[781] = inter_3[781];
    assign inter_4[782] = inter_3[782];
    assign inter_4[783] = inter_3[783];
    assign inter_4[784] = inter_3[784]^inter_3[792];
    assign inter_4[785] = inter_3[785]^inter_3[793];
    assign inter_4[786] = inter_3[786]^inter_3[794];
    assign inter_4[787] = inter_3[787]^inter_3[795];
    assign inter_4[788] = inter_3[788]^inter_3[796];
    assign inter_4[789] = inter_3[789]^inter_3[797];
    assign inter_4[790] = inter_3[790]^inter_3[798];
    assign inter_4[791] = inter_3[791]^inter_3[799];
    assign inter_4[792] = inter_3[792];
    assign inter_4[793] = inter_3[793];
    assign inter_4[794] = inter_3[794];
    assign inter_4[795] = inter_3[795];
    assign inter_4[796] = inter_3[796];
    assign inter_4[797] = inter_3[797];
    assign inter_4[798] = inter_3[798];
    assign inter_4[799] = inter_3[799];
    assign inter_4[800] = inter_3[800]^inter_3[808];
    assign inter_4[801] = inter_3[801]^inter_3[809];
    assign inter_4[802] = inter_3[802]^inter_3[810];
    assign inter_4[803] = inter_3[803]^inter_3[811];
    assign inter_4[804] = inter_3[804]^inter_3[812];
    assign inter_4[805] = inter_3[805]^inter_3[813];
    assign inter_4[806] = inter_3[806]^inter_3[814];
    assign inter_4[807] = inter_3[807]^inter_3[815];
    assign inter_4[808] = inter_3[808];
    assign inter_4[809] = inter_3[809];
    assign inter_4[810] = inter_3[810];
    assign inter_4[811] = inter_3[811];
    assign inter_4[812] = inter_3[812];
    assign inter_4[813] = inter_3[813];
    assign inter_4[814] = inter_3[814];
    assign inter_4[815] = inter_3[815];
    assign inter_4[816] = inter_3[816]^inter_3[824];
    assign inter_4[817] = inter_3[817]^inter_3[825];
    assign inter_4[818] = inter_3[818]^inter_3[826];
    assign inter_4[819] = inter_3[819]^inter_3[827];
    assign inter_4[820] = inter_3[820]^inter_3[828];
    assign inter_4[821] = inter_3[821]^inter_3[829];
    assign inter_4[822] = inter_3[822]^inter_3[830];
    assign inter_4[823] = inter_3[823]^inter_3[831];
    assign inter_4[824] = inter_3[824];
    assign inter_4[825] = inter_3[825];
    assign inter_4[826] = inter_3[826];
    assign inter_4[827] = inter_3[827];
    assign inter_4[828] = inter_3[828];
    assign inter_4[829] = inter_3[829];
    assign inter_4[830] = inter_3[830];
    assign inter_4[831] = inter_3[831];
    assign inter_4[832] = inter_3[832]^inter_3[840];
    assign inter_4[833] = inter_3[833]^inter_3[841];
    assign inter_4[834] = inter_3[834]^inter_3[842];
    assign inter_4[835] = inter_3[835]^inter_3[843];
    assign inter_4[836] = inter_3[836]^inter_3[844];
    assign inter_4[837] = inter_3[837]^inter_3[845];
    assign inter_4[838] = inter_3[838]^inter_3[846];
    assign inter_4[839] = inter_3[839]^inter_3[847];
    assign inter_4[840] = inter_3[840];
    assign inter_4[841] = inter_3[841];
    assign inter_4[842] = inter_3[842];
    assign inter_4[843] = inter_3[843];
    assign inter_4[844] = inter_3[844];
    assign inter_4[845] = inter_3[845];
    assign inter_4[846] = inter_3[846];
    assign inter_4[847] = inter_3[847];
    assign inter_4[848] = inter_3[848]^inter_3[856];
    assign inter_4[849] = inter_3[849]^inter_3[857];
    assign inter_4[850] = inter_3[850]^inter_3[858];
    assign inter_4[851] = inter_3[851]^inter_3[859];
    assign inter_4[852] = inter_3[852]^inter_3[860];
    assign inter_4[853] = inter_3[853]^inter_3[861];
    assign inter_4[854] = inter_3[854]^inter_3[862];
    assign inter_4[855] = inter_3[855]^inter_3[863];
    assign inter_4[856] = inter_3[856];
    assign inter_4[857] = inter_3[857];
    assign inter_4[858] = inter_3[858];
    assign inter_4[859] = inter_3[859];
    assign inter_4[860] = inter_3[860];
    assign inter_4[861] = inter_3[861];
    assign inter_4[862] = inter_3[862];
    assign inter_4[863] = inter_3[863];
    assign inter_4[864] = inter_3[864]^inter_3[872];
    assign inter_4[865] = inter_3[865]^inter_3[873];
    assign inter_4[866] = inter_3[866]^inter_3[874];
    assign inter_4[867] = inter_3[867]^inter_3[875];
    assign inter_4[868] = inter_3[868]^inter_3[876];
    assign inter_4[869] = inter_3[869]^inter_3[877];
    assign inter_4[870] = inter_3[870]^inter_3[878];
    assign inter_4[871] = inter_3[871]^inter_3[879];
    assign inter_4[872] = inter_3[872];
    assign inter_4[873] = inter_3[873];
    assign inter_4[874] = inter_3[874];
    assign inter_4[875] = inter_3[875];
    assign inter_4[876] = inter_3[876];
    assign inter_4[877] = inter_3[877];
    assign inter_4[878] = inter_3[878];
    assign inter_4[879] = inter_3[879];
    assign inter_4[880] = inter_3[880]^inter_3[888];
    assign inter_4[881] = inter_3[881]^inter_3[889];
    assign inter_4[882] = inter_3[882]^inter_3[890];
    assign inter_4[883] = inter_3[883]^inter_3[891];
    assign inter_4[884] = inter_3[884]^inter_3[892];
    assign inter_4[885] = inter_3[885]^inter_3[893];
    assign inter_4[886] = inter_3[886]^inter_3[894];
    assign inter_4[887] = inter_3[887]^inter_3[895];
    assign inter_4[888] = inter_3[888];
    assign inter_4[889] = inter_3[889];
    assign inter_4[890] = inter_3[890];
    assign inter_4[891] = inter_3[891];
    assign inter_4[892] = inter_3[892];
    assign inter_4[893] = inter_3[893];
    assign inter_4[894] = inter_3[894];
    assign inter_4[895] = inter_3[895];
    assign inter_4[896] = inter_3[896]^inter_3[904];
    assign inter_4[897] = inter_3[897]^inter_3[905];
    assign inter_4[898] = inter_3[898]^inter_3[906];
    assign inter_4[899] = inter_3[899]^inter_3[907];
    assign inter_4[900] = inter_3[900]^inter_3[908];
    assign inter_4[901] = inter_3[901]^inter_3[909];
    assign inter_4[902] = inter_3[902]^inter_3[910];
    assign inter_4[903] = inter_3[903]^inter_3[911];
    assign inter_4[904] = inter_3[904];
    assign inter_4[905] = inter_3[905];
    assign inter_4[906] = inter_3[906];
    assign inter_4[907] = inter_3[907];
    assign inter_4[908] = inter_3[908];
    assign inter_4[909] = inter_3[909];
    assign inter_4[910] = inter_3[910];
    assign inter_4[911] = inter_3[911];
    assign inter_4[912] = inter_3[912]^inter_3[920];
    assign inter_4[913] = inter_3[913]^inter_3[921];
    assign inter_4[914] = inter_3[914]^inter_3[922];
    assign inter_4[915] = inter_3[915]^inter_3[923];
    assign inter_4[916] = inter_3[916]^inter_3[924];
    assign inter_4[917] = inter_3[917]^inter_3[925];
    assign inter_4[918] = inter_3[918]^inter_3[926];
    assign inter_4[919] = inter_3[919]^inter_3[927];
    assign inter_4[920] = inter_3[920];
    assign inter_4[921] = inter_3[921];
    assign inter_4[922] = inter_3[922];
    assign inter_4[923] = inter_3[923];
    assign inter_4[924] = inter_3[924];
    assign inter_4[925] = inter_3[925];
    assign inter_4[926] = inter_3[926];
    assign inter_4[927] = inter_3[927];
    assign inter_4[928] = inter_3[928]^inter_3[936];
    assign inter_4[929] = inter_3[929]^inter_3[937];
    assign inter_4[930] = inter_3[930]^inter_3[938];
    assign inter_4[931] = inter_3[931]^inter_3[939];
    assign inter_4[932] = inter_3[932]^inter_3[940];
    assign inter_4[933] = inter_3[933]^inter_3[941];
    assign inter_4[934] = inter_3[934]^inter_3[942];
    assign inter_4[935] = inter_3[935]^inter_3[943];
    assign inter_4[936] = inter_3[936];
    assign inter_4[937] = inter_3[937];
    assign inter_4[938] = inter_3[938];
    assign inter_4[939] = inter_3[939];
    assign inter_4[940] = inter_3[940];
    assign inter_4[941] = inter_3[941];
    assign inter_4[942] = inter_3[942];
    assign inter_4[943] = inter_3[943];
    assign inter_4[944] = inter_3[944]^inter_3[952];
    assign inter_4[945] = inter_3[945]^inter_3[953];
    assign inter_4[946] = inter_3[946]^inter_3[954];
    assign inter_4[947] = inter_3[947]^inter_3[955];
    assign inter_4[948] = inter_3[948]^inter_3[956];
    assign inter_4[949] = inter_3[949]^inter_3[957];
    assign inter_4[950] = inter_3[950]^inter_3[958];
    assign inter_4[951] = inter_3[951]^inter_3[959];
    assign inter_4[952] = inter_3[952];
    assign inter_4[953] = inter_3[953];
    assign inter_4[954] = inter_3[954];
    assign inter_4[955] = inter_3[955];
    assign inter_4[956] = inter_3[956];
    assign inter_4[957] = inter_3[957];
    assign inter_4[958] = inter_3[958];
    assign inter_4[959] = inter_3[959];
    assign inter_4[960] = inter_3[960]^inter_3[968];
    assign inter_4[961] = inter_3[961]^inter_3[969];
    assign inter_4[962] = inter_3[962]^inter_3[970];
    assign inter_4[963] = inter_3[963]^inter_3[971];
    assign inter_4[964] = inter_3[964]^inter_3[972];
    assign inter_4[965] = inter_3[965]^inter_3[973];
    assign inter_4[966] = inter_3[966]^inter_3[974];
    assign inter_4[967] = inter_3[967]^inter_3[975];
    assign inter_4[968] = inter_3[968];
    assign inter_4[969] = inter_3[969];
    assign inter_4[970] = inter_3[970];
    assign inter_4[971] = inter_3[971];
    assign inter_4[972] = inter_3[972];
    assign inter_4[973] = inter_3[973];
    assign inter_4[974] = inter_3[974];
    assign inter_4[975] = inter_3[975];
    assign inter_4[976] = inter_3[976]^inter_3[984];
    assign inter_4[977] = inter_3[977]^inter_3[985];
    assign inter_4[978] = inter_3[978]^inter_3[986];
    assign inter_4[979] = inter_3[979]^inter_3[987];
    assign inter_4[980] = inter_3[980]^inter_3[988];
    assign inter_4[981] = inter_3[981]^inter_3[989];
    assign inter_4[982] = inter_3[982]^inter_3[990];
    assign inter_4[983] = inter_3[983]^inter_3[991];
    assign inter_4[984] = inter_3[984];
    assign inter_4[985] = inter_3[985];
    assign inter_4[986] = inter_3[986];
    assign inter_4[987] = inter_3[987];
    assign inter_4[988] = inter_3[988];
    assign inter_4[989] = inter_3[989];
    assign inter_4[990] = inter_3[990];
    assign inter_4[991] = inter_3[991];
    assign inter_4[992] = inter_3[992]^inter_3[1000];
    assign inter_4[993] = inter_3[993]^inter_3[1001];
    assign inter_4[994] = inter_3[994]^inter_3[1002];
    assign inter_4[995] = inter_3[995]^inter_3[1003];
    assign inter_4[996] = inter_3[996]^inter_3[1004];
    assign inter_4[997] = inter_3[997]^inter_3[1005];
    assign inter_4[998] = inter_3[998]^inter_3[1006];
    assign inter_4[999] = inter_3[999]^inter_3[1007];
    assign inter_4[1000] = inter_3[1000];
    assign inter_4[1001] = inter_3[1001];
    assign inter_4[1002] = inter_3[1002];
    assign inter_4[1003] = inter_3[1003];
    assign inter_4[1004] = inter_3[1004];
    assign inter_4[1005] = inter_3[1005];
    assign inter_4[1006] = inter_3[1006];
    assign inter_4[1007] = inter_3[1007];
    assign inter_4[1008] = inter_3[1008]^inter_3[1016];
    assign inter_4[1009] = inter_3[1009]^inter_3[1017];
    assign inter_4[1010] = inter_3[1010]^inter_3[1018];
    assign inter_4[1011] = inter_3[1011]^inter_3[1019];
    assign inter_4[1012] = inter_3[1012]^inter_3[1020];
    assign inter_4[1013] = inter_3[1013]^inter_3[1021];
    assign inter_4[1014] = inter_3[1014]^inter_3[1022];
    assign inter_4[1015] = inter_3[1015]^inter_3[1023];
    assign inter_4[1016] = inter_3[1016];
    assign inter_4[1017] = inter_3[1017];
    assign inter_4[1018] = inter_3[1018];
    assign inter_4[1019] = inter_3[1019];
    assign inter_4[1020] = inter_3[1020];
    assign inter_4[1021] = inter_3[1021];
    assign inter_4[1022] = inter_3[1022];
    assign inter_4[1023] = inter_3[1023];
    /***************************/
    assign inter_5[0] = inter_4[0]^inter_4[16];
    assign inter_5[1] = inter_4[1]^inter_4[17];
    assign inter_5[2] = inter_4[2]^inter_4[18];
    assign inter_5[3] = inter_4[3]^inter_4[19];
    assign inter_5[4] = inter_4[4]^inter_4[20];
    assign inter_5[5] = inter_4[5]^inter_4[21];
    assign inter_5[6] = inter_4[6]^inter_4[22];
    assign inter_5[7] = inter_4[7]^inter_4[23];
    assign inter_5[8] = inter_4[8]^inter_4[24];
    assign inter_5[9] = inter_4[9]^inter_4[25];
    assign inter_5[10] = inter_4[10]^inter_4[26];
    assign inter_5[11] = inter_4[11]^inter_4[27];
    assign inter_5[12] = inter_4[12]^inter_4[28];
    assign inter_5[13] = inter_4[13]^inter_4[29];
    assign inter_5[14] = inter_4[14]^inter_4[30];
    assign inter_5[15] = inter_4[15]^inter_4[31];
    assign inter_5[16] = inter_4[16];
    assign inter_5[17] = inter_4[17];
    assign inter_5[18] = inter_4[18];
    assign inter_5[19] = inter_4[19];
    assign inter_5[20] = inter_4[20];
    assign inter_5[21] = inter_4[21];
    assign inter_5[22] = inter_4[22];
    assign inter_5[23] = inter_4[23];
    assign inter_5[24] = inter_4[24];
    assign inter_5[25] = inter_4[25];
    assign inter_5[26] = inter_4[26];
    assign inter_5[27] = inter_4[27];
    assign inter_5[28] = inter_4[28];
    assign inter_5[29] = inter_4[29];
    assign inter_5[30] = inter_4[30];
    assign inter_5[31] = inter_4[31];
    assign inter_5[32] = inter_4[32]^inter_4[48];
    assign inter_5[33] = inter_4[33]^inter_4[49];
    assign inter_5[34] = inter_4[34]^inter_4[50];
    assign inter_5[35] = inter_4[35]^inter_4[51];
    assign inter_5[36] = inter_4[36]^inter_4[52];
    assign inter_5[37] = inter_4[37]^inter_4[53];
    assign inter_5[38] = inter_4[38]^inter_4[54];
    assign inter_5[39] = inter_4[39]^inter_4[55];
    assign inter_5[40] = inter_4[40]^inter_4[56];
    assign inter_5[41] = inter_4[41]^inter_4[57];
    assign inter_5[42] = inter_4[42]^inter_4[58];
    assign inter_5[43] = inter_4[43]^inter_4[59];
    assign inter_5[44] = inter_4[44]^inter_4[60];
    assign inter_5[45] = inter_4[45]^inter_4[61];
    assign inter_5[46] = inter_4[46]^inter_4[62];
    assign inter_5[47] = inter_4[47]^inter_4[63];
    assign inter_5[48] = inter_4[48];
    assign inter_5[49] = inter_4[49];
    assign inter_5[50] = inter_4[50];
    assign inter_5[51] = inter_4[51];
    assign inter_5[52] = inter_4[52];
    assign inter_5[53] = inter_4[53];
    assign inter_5[54] = inter_4[54];
    assign inter_5[55] = inter_4[55];
    assign inter_5[56] = inter_4[56];
    assign inter_5[57] = inter_4[57];
    assign inter_5[58] = inter_4[58];
    assign inter_5[59] = inter_4[59];
    assign inter_5[60] = inter_4[60];
    assign inter_5[61] = inter_4[61];
    assign inter_5[62] = inter_4[62];
    assign inter_5[63] = inter_4[63];
    assign inter_5[64] = inter_4[64]^inter_4[80];
    assign inter_5[65] = inter_4[65]^inter_4[81];
    assign inter_5[66] = inter_4[66]^inter_4[82];
    assign inter_5[67] = inter_4[67]^inter_4[83];
    assign inter_5[68] = inter_4[68]^inter_4[84];
    assign inter_5[69] = inter_4[69]^inter_4[85];
    assign inter_5[70] = inter_4[70]^inter_4[86];
    assign inter_5[71] = inter_4[71]^inter_4[87];
    assign inter_5[72] = inter_4[72]^inter_4[88];
    assign inter_5[73] = inter_4[73]^inter_4[89];
    assign inter_5[74] = inter_4[74]^inter_4[90];
    assign inter_5[75] = inter_4[75]^inter_4[91];
    assign inter_5[76] = inter_4[76]^inter_4[92];
    assign inter_5[77] = inter_4[77]^inter_4[93];
    assign inter_5[78] = inter_4[78]^inter_4[94];
    assign inter_5[79] = inter_4[79]^inter_4[95];
    assign inter_5[80] = inter_4[80];
    assign inter_5[81] = inter_4[81];
    assign inter_5[82] = inter_4[82];
    assign inter_5[83] = inter_4[83];
    assign inter_5[84] = inter_4[84];
    assign inter_5[85] = inter_4[85];
    assign inter_5[86] = inter_4[86];
    assign inter_5[87] = inter_4[87];
    assign inter_5[88] = inter_4[88];
    assign inter_5[89] = inter_4[89];
    assign inter_5[90] = inter_4[90];
    assign inter_5[91] = inter_4[91];
    assign inter_5[92] = inter_4[92];
    assign inter_5[93] = inter_4[93];
    assign inter_5[94] = inter_4[94];
    assign inter_5[95] = inter_4[95];
    assign inter_5[96] = inter_4[96]^inter_4[112];
    assign inter_5[97] = inter_4[97]^inter_4[113];
    assign inter_5[98] = inter_4[98]^inter_4[114];
    assign inter_5[99] = inter_4[99]^inter_4[115];
    assign inter_5[100] = inter_4[100]^inter_4[116];
    assign inter_5[101] = inter_4[101]^inter_4[117];
    assign inter_5[102] = inter_4[102]^inter_4[118];
    assign inter_5[103] = inter_4[103]^inter_4[119];
    assign inter_5[104] = inter_4[104]^inter_4[120];
    assign inter_5[105] = inter_4[105]^inter_4[121];
    assign inter_5[106] = inter_4[106]^inter_4[122];
    assign inter_5[107] = inter_4[107]^inter_4[123];
    assign inter_5[108] = inter_4[108]^inter_4[124];
    assign inter_5[109] = inter_4[109]^inter_4[125];
    assign inter_5[110] = inter_4[110]^inter_4[126];
    assign inter_5[111] = inter_4[111]^inter_4[127];
    assign inter_5[112] = inter_4[112];
    assign inter_5[113] = inter_4[113];
    assign inter_5[114] = inter_4[114];
    assign inter_5[115] = inter_4[115];
    assign inter_5[116] = inter_4[116];
    assign inter_5[117] = inter_4[117];
    assign inter_5[118] = inter_4[118];
    assign inter_5[119] = inter_4[119];
    assign inter_5[120] = inter_4[120];
    assign inter_5[121] = inter_4[121];
    assign inter_5[122] = inter_4[122];
    assign inter_5[123] = inter_4[123];
    assign inter_5[124] = inter_4[124];
    assign inter_5[125] = inter_4[125];
    assign inter_5[126] = inter_4[126];
    assign inter_5[127] = inter_4[127];
    assign inter_5[128] = inter_4[128]^inter_4[144];
    assign inter_5[129] = inter_4[129]^inter_4[145];
    assign inter_5[130] = inter_4[130]^inter_4[146];
    assign inter_5[131] = inter_4[131]^inter_4[147];
    assign inter_5[132] = inter_4[132]^inter_4[148];
    assign inter_5[133] = inter_4[133]^inter_4[149];
    assign inter_5[134] = inter_4[134]^inter_4[150];
    assign inter_5[135] = inter_4[135]^inter_4[151];
    assign inter_5[136] = inter_4[136]^inter_4[152];
    assign inter_5[137] = inter_4[137]^inter_4[153];
    assign inter_5[138] = inter_4[138]^inter_4[154];
    assign inter_5[139] = inter_4[139]^inter_4[155];
    assign inter_5[140] = inter_4[140]^inter_4[156];
    assign inter_5[141] = inter_4[141]^inter_4[157];
    assign inter_5[142] = inter_4[142]^inter_4[158];
    assign inter_5[143] = inter_4[143]^inter_4[159];
    assign inter_5[144] = inter_4[144];
    assign inter_5[145] = inter_4[145];
    assign inter_5[146] = inter_4[146];
    assign inter_5[147] = inter_4[147];
    assign inter_5[148] = inter_4[148];
    assign inter_5[149] = inter_4[149];
    assign inter_5[150] = inter_4[150];
    assign inter_5[151] = inter_4[151];
    assign inter_5[152] = inter_4[152];
    assign inter_5[153] = inter_4[153];
    assign inter_5[154] = inter_4[154];
    assign inter_5[155] = inter_4[155];
    assign inter_5[156] = inter_4[156];
    assign inter_5[157] = inter_4[157];
    assign inter_5[158] = inter_4[158];
    assign inter_5[159] = inter_4[159];
    assign inter_5[160] = inter_4[160]^inter_4[176];
    assign inter_5[161] = inter_4[161]^inter_4[177];
    assign inter_5[162] = inter_4[162]^inter_4[178];
    assign inter_5[163] = inter_4[163]^inter_4[179];
    assign inter_5[164] = inter_4[164]^inter_4[180];
    assign inter_5[165] = inter_4[165]^inter_4[181];
    assign inter_5[166] = inter_4[166]^inter_4[182];
    assign inter_5[167] = inter_4[167]^inter_4[183];
    assign inter_5[168] = inter_4[168]^inter_4[184];
    assign inter_5[169] = inter_4[169]^inter_4[185];
    assign inter_5[170] = inter_4[170]^inter_4[186];
    assign inter_5[171] = inter_4[171]^inter_4[187];
    assign inter_5[172] = inter_4[172]^inter_4[188];
    assign inter_5[173] = inter_4[173]^inter_4[189];
    assign inter_5[174] = inter_4[174]^inter_4[190];
    assign inter_5[175] = inter_4[175]^inter_4[191];
    assign inter_5[176] = inter_4[176];
    assign inter_5[177] = inter_4[177];
    assign inter_5[178] = inter_4[178];
    assign inter_5[179] = inter_4[179];
    assign inter_5[180] = inter_4[180];
    assign inter_5[181] = inter_4[181];
    assign inter_5[182] = inter_4[182];
    assign inter_5[183] = inter_4[183];
    assign inter_5[184] = inter_4[184];
    assign inter_5[185] = inter_4[185];
    assign inter_5[186] = inter_4[186];
    assign inter_5[187] = inter_4[187];
    assign inter_5[188] = inter_4[188];
    assign inter_5[189] = inter_4[189];
    assign inter_5[190] = inter_4[190];
    assign inter_5[191] = inter_4[191];
    assign inter_5[192] = inter_4[192]^inter_4[208];
    assign inter_5[193] = inter_4[193]^inter_4[209];
    assign inter_5[194] = inter_4[194]^inter_4[210];
    assign inter_5[195] = inter_4[195]^inter_4[211];
    assign inter_5[196] = inter_4[196]^inter_4[212];
    assign inter_5[197] = inter_4[197]^inter_4[213];
    assign inter_5[198] = inter_4[198]^inter_4[214];
    assign inter_5[199] = inter_4[199]^inter_4[215];
    assign inter_5[200] = inter_4[200]^inter_4[216];
    assign inter_5[201] = inter_4[201]^inter_4[217];
    assign inter_5[202] = inter_4[202]^inter_4[218];
    assign inter_5[203] = inter_4[203]^inter_4[219];
    assign inter_5[204] = inter_4[204]^inter_4[220];
    assign inter_5[205] = inter_4[205]^inter_4[221];
    assign inter_5[206] = inter_4[206]^inter_4[222];
    assign inter_5[207] = inter_4[207]^inter_4[223];
    assign inter_5[208] = inter_4[208];
    assign inter_5[209] = inter_4[209];
    assign inter_5[210] = inter_4[210];
    assign inter_5[211] = inter_4[211];
    assign inter_5[212] = inter_4[212];
    assign inter_5[213] = inter_4[213];
    assign inter_5[214] = inter_4[214];
    assign inter_5[215] = inter_4[215];
    assign inter_5[216] = inter_4[216];
    assign inter_5[217] = inter_4[217];
    assign inter_5[218] = inter_4[218];
    assign inter_5[219] = inter_4[219];
    assign inter_5[220] = inter_4[220];
    assign inter_5[221] = inter_4[221];
    assign inter_5[222] = inter_4[222];
    assign inter_5[223] = inter_4[223];
    assign inter_5[224] = inter_4[224]^inter_4[240];
    assign inter_5[225] = inter_4[225]^inter_4[241];
    assign inter_5[226] = inter_4[226]^inter_4[242];
    assign inter_5[227] = inter_4[227]^inter_4[243];
    assign inter_5[228] = inter_4[228]^inter_4[244];
    assign inter_5[229] = inter_4[229]^inter_4[245];
    assign inter_5[230] = inter_4[230]^inter_4[246];
    assign inter_5[231] = inter_4[231]^inter_4[247];
    assign inter_5[232] = inter_4[232]^inter_4[248];
    assign inter_5[233] = inter_4[233]^inter_4[249];
    assign inter_5[234] = inter_4[234]^inter_4[250];
    assign inter_5[235] = inter_4[235]^inter_4[251];
    assign inter_5[236] = inter_4[236]^inter_4[252];
    assign inter_5[237] = inter_4[237]^inter_4[253];
    assign inter_5[238] = inter_4[238]^inter_4[254];
    assign inter_5[239] = inter_4[239]^inter_4[255];
    assign inter_5[240] = inter_4[240];
    assign inter_5[241] = inter_4[241];
    assign inter_5[242] = inter_4[242];
    assign inter_5[243] = inter_4[243];
    assign inter_5[244] = inter_4[244];
    assign inter_5[245] = inter_4[245];
    assign inter_5[246] = inter_4[246];
    assign inter_5[247] = inter_4[247];
    assign inter_5[248] = inter_4[248];
    assign inter_5[249] = inter_4[249];
    assign inter_5[250] = inter_4[250];
    assign inter_5[251] = inter_4[251];
    assign inter_5[252] = inter_4[252];
    assign inter_5[253] = inter_4[253];
    assign inter_5[254] = inter_4[254];
    assign inter_5[255] = inter_4[255];
    assign inter_5[256] = inter_4[256]^inter_4[272];
    assign inter_5[257] = inter_4[257]^inter_4[273];
    assign inter_5[258] = inter_4[258]^inter_4[274];
    assign inter_5[259] = inter_4[259]^inter_4[275];
    assign inter_5[260] = inter_4[260]^inter_4[276];
    assign inter_5[261] = inter_4[261]^inter_4[277];
    assign inter_5[262] = inter_4[262]^inter_4[278];
    assign inter_5[263] = inter_4[263]^inter_4[279];
    assign inter_5[264] = inter_4[264]^inter_4[280];
    assign inter_5[265] = inter_4[265]^inter_4[281];
    assign inter_5[266] = inter_4[266]^inter_4[282];
    assign inter_5[267] = inter_4[267]^inter_4[283];
    assign inter_5[268] = inter_4[268]^inter_4[284];
    assign inter_5[269] = inter_4[269]^inter_4[285];
    assign inter_5[270] = inter_4[270]^inter_4[286];
    assign inter_5[271] = inter_4[271]^inter_4[287];
    assign inter_5[272] = inter_4[272];
    assign inter_5[273] = inter_4[273];
    assign inter_5[274] = inter_4[274];
    assign inter_5[275] = inter_4[275];
    assign inter_5[276] = inter_4[276];
    assign inter_5[277] = inter_4[277];
    assign inter_5[278] = inter_4[278];
    assign inter_5[279] = inter_4[279];
    assign inter_5[280] = inter_4[280];
    assign inter_5[281] = inter_4[281];
    assign inter_5[282] = inter_4[282];
    assign inter_5[283] = inter_4[283];
    assign inter_5[284] = inter_4[284];
    assign inter_5[285] = inter_4[285];
    assign inter_5[286] = inter_4[286];
    assign inter_5[287] = inter_4[287];
    assign inter_5[288] = inter_4[288]^inter_4[304];
    assign inter_5[289] = inter_4[289]^inter_4[305];
    assign inter_5[290] = inter_4[290]^inter_4[306];
    assign inter_5[291] = inter_4[291]^inter_4[307];
    assign inter_5[292] = inter_4[292]^inter_4[308];
    assign inter_5[293] = inter_4[293]^inter_4[309];
    assign inter_5[294] = inter_4[294]^inter_4[310];
    assign inter_5[295] = inter_4[295]^inter_4[311];
    assign inter_5[296] = inter_4[296]^inter_4[312];
    assign inter_5[297] = inter_4[297]^inter_4[313];
    assign inter_5[298] = inter_4[298]^inter_4[314];
    assign inter_5[299] = inter_4[299]^inter_4[315];
    assign inter_5[300] = inter_4[300]^inter_4[316];
    assign inter_5[301] = inter_4[301]^inter_4[317];
    assign inter_5[302] = inter_4[302]^inter_4[318];
    assign inter_5[303] = inter_4[303]^inter_4[319];
    assign inter_5[304] = inter_4[304];
    assign inter_5[305] = inter_4[305];
    assign inter_5[306] = inter_4[306];
    assign inter_5[307] = inter_4[307];
    assign inter_5[308] = inter_4[308];
    assign inter_5[309] = inter_4[309];
    assign inter_5[310] = inter_4[310];
    assign inter_5[311] = inter_4[311];
    assign inter_5[312] = inter_4[312];
    assign inter_5[313] = inter_4[313];
    assign inter_5[314] = inter_4[314];
    assign inter_5[315] = inter_4[315];
    assign inter_5[316] = inter_4[316];
    assign inter_5[317] = inter_4[317];
    assign inter_5[318] = inter_4[318];
    assign inter_5[319] = inter_4[319];
    assign inter_5[320] = inter_4[320]^inter_4[336];
    assign inter_5[321] = inter_4[321]^inter_4[337];
    assign inter_5[322] = inter_4[322]^inter_4[338];
    assign inter_5[323] = inter_4[323]^inter_4[339];
    assign inter_5[324] = inter_4[324]^inter_4[340];
    assign inter_5[325] = inter_4[325]^inter_4[341];
    assign inter_5[326] = inter_4[326]^inter_4[342];
    assign inter_5[327] = inter_4[327]^inter_4[343];
    assign inter_5[328] = inter_4[328]^inter_4[344];
    assign inter_5[329] = inter_4[329]^inter_4[345];
    assign inter_5[330] = inter_4[330]^inter_4[346];
    assign inter_5[331] = inter_4[331]^inter_4[347];
    assign inter_5[332] = inter_4[332]^inter_4[348];
    assign inter_5[333] = inter_4[333]^inter_4[349];
    assign inter_5[334] = inter_4[334]^inter_4[350];
    assign inter_5[335] = inter_4[335]^inter_4[351];
    assign inter_5[336] = inter_4[336];
    assign inter_5[337] = inter_4[337];
    assign inter_5[338] = inter_4[338];
    assign inter_5[339] = inter_4[339];
    assign inter_5[340] = inter_4[340];
    assign inter_5[341] = inter_4[341];
    assign inter_5[342] = inter_4[342];
    assign inter_5[343] = inter_4[343];
    assign inter_5[344] = inter_4[344];
    assign inter_5[345] = inter_4[345];
    assign inter_5[346] = inter_4[346];
    assign inter_5[347] = inter_4[347];
    assign inter_5[348] = inter_4[348];
    assign inter_5[349] = inter_4[349];
    assign inter_5[350] = inter_4[350];
    assign inter_5[351] = inter_4[351];
    assign inter_5[352] = inter_4[352]^inter_4[368];
    assign inter_5[353] = inter_4[353]^inter_4[369];
    assign inter_5[354] = inter_4[354]^inter_4[370];
    assign inter_5[355] = inter_4[355]^inter_4[371];
    assign inter_5[356] = inter_4[356]^inter_4[372];
    assign inter_5[357] = inter_4[357]^inter_4[373];
    assign inter_5[358] = inter_4[358]^inter_4[374];
    assign inter_5[359] = inter_4[359]^inter_4[375];
    assign inter_5[360] = inter_4[360]^inter_4[376];
    assign inter_5[361] = inter_4[361]^inter_4[377];
    assign inter_5[362] = inter_4[362]^inter_4[378];
    assign inter_5[363] = inter_4[363]^inter_4[379];
    assign inter_5[364] = inter_4[364]^inter_4[380];
    assign inter_5[365] = inter_4[365]^inter_4[381];
    assign inter_5[366] = inter_4[366]^inter_4[382];
    assign inter_5[367] = inter_4[367]^inter_4[383];
    assign inter_5[368] = inter_4[368];
    assign inter_5[369] = inter_4[369];
    assign inter_5[370] = inter_4[370];
    assign inter_5[371] = inter_4[371];
    assign inter_5[372] = inter_4[372];
    assign inter_5[373] = inter_4[373];
    assign inter_5[374] = inter_4[374];
    assign inter_5[375] = inter_4[375];
    assign inter_5[376] = inter_4[376];
    assign inter_5[377] = inter_4[377];
    assign inter_5[378] = inter_4[378];
    assign inter_5[379] = inter_4[379];
    assign inter_5[380] = inter_4[380];
    assign inter_5[381] = inter_4[381];
    assign inter_5[382] = inter_4[382];
    assign inter_5[383] = inter_4[383];
    assign inter_5[384] = inter_4[384]^inter_4[400];
    assign inter_5[385] = inter_4[385]^inter_4[401];
    assign inter_5[386] = inter_4[386]^inter_4[402];
    assign inter_5[387] = inter_4[387]^inter_4[403];
    assign inter_5[388] = inter_4[388]^inter_4[404];
    assign inter_5[389] = inter_4[389]^inter_4[405];
    assign inter_5[390] = inter_4[390]^inter_4[406];
    assign inter_5[391] = inter_4[391]^inter_4[407];
    assign inter_5[392] = inter_4[392]^inter_4[408];
    assign inter_5[393] = inter_4[393]^inter_4[409];
    assign inter_5[394] = inter_4[394]^inter_4[410];
    assign inter_5[395] = inter_4[395]^inter_4[411];
    assign inter_5[396] = inter_4[396]^inter_4[412];
    assign inter_5[397] = inter_4[397]^inter_4[413];
    assign inter_5[398] = inter_4[398]^inter_4[414];
    assign inter_5[399] = inter_4[399]^inter_4[415];
    assign inter_5[400] = inter_4[400];
    assign inter_5[401] = inter_4[401];
    assign inter_5[402] = inter_4[402];
    assign inter_5[403] = inter_4[403];
    assign inter_5[404] = inter_4[404];
    assign inter_5[405] = inter_4[405];
    assign inter_5[406] = inter_4[406];
    assign inter_5[407] = inter_4[407];
    assign inter_5[408] = inter_4[408];
    assign inter_5[409] = inter_4[409];
    assign inter_5[410] = inter_4[410];
    assign inter_5[411] = inter_4[411];
    assign inter_5[412] = inter_4[412];
    assign inter_5[413] = inter_4[413];
    assign inter_5[414] = inter_4[414];
    assign inter_5[415] = inter_4[415];
    assign inter_5[416] = inter_4[416]^inter_4[432];
    assign inter_5[417] = inter_4[417]^inter_4[433];
    assign inter_5[418] = inter_4[418]^inter_4[434];
    assign inter_5[419] = inter_4[419]^inter_4[435];
    assign inter_5[420] = inter_4[420]^inter_4[436];
    assign inter_5[421] = inter_4[421]^inter_4[437];
    assign inter_5[422] = inter_4[422]^inter_4[438];
    assign inter_5[423] = inter_4[423]^inter_4[439];
    assign inter_5[424] = inter_4[424]^inter_4[440];
    assign inter_5[425] = inter_4[425]^inter_4[441];
    assign inter_5[426] = inter_4[426]^inter_4[442];
    assign inter_5[427] = inter_4[427]^inter_4[443];
    assign inter_5[428] = inter_4[428]^inter_4[444];
    assign inter_5[429] = inter_4[429]^inter_4[445];
    assign inter_5[430] = inter_4[430]^inter_4[446];
    assign inter_5[431] = inter_4[431]^inter_4[447];
    assign inter_5[432] = inter_4[432];
    assign inter_5[433] = inter_4[433];
    assign inter_5[434] = inter_4[434];
    assign inter_5[435] = inter_4[435];
    assign inter_5[436] = inter_4[436];
    assign inter_5[437] = inter_4[437];
    assign inter_5[438] = inter_4[438];
    assign inter_5[439] = inter_4[439];
    assign inter_5[440] = inter_4[440];
    assign inter_5[441] = inter_4[441];
    assign inter_5[442] = inter_4[442];
    assign inter_5[443] = inter_4[443];
    assign inter_5[444] = inter_4[444];
    assign inter_5[445] = inter_4[445];
    assign inter_5[446] = inter_4[446];
    assign inter_5[447] = inter_4[447];
    assign inter_5[448] = inter_4[448]^inter_4[464];
    assign inter_5[449] = inter_4[449]^inter_4[465];
    assign inter_5[450] = inter_4[450]^inter_4[466];
    assign inter_5[451] = inter_4[451]^inter_4[467];
    assign inter_5[452] = inter_4[452]^inter_4[468];
    assign inter_5[453] = inter_4[453]^inter_4[469];
    assign inter_5[454] = inter_4[454]^inter_4[470];
    assign inter_5[455] = inter_4[455]^inter_4[471];
    assign inter_5[456] = inter_4[456]^inter_4[472];
    assign inter_5[457] = inter_4[457]^inter_4[473];
    assign inter_5[458] = inter_4[458]^inter_4[474];
    assign inter_5[459] = inter_4[459]^inter_4[475];
    assign inter_5[460] = inter_4[460]^inter_4[476];
    assign inter_5[461] = inter_4[461]^inter_4[477];
    assign inter_5[462] = inter_4[462]^inter_4[478];
    assign inter_5[463] = inter_4[463]^inter_4[479];
    assign inter_5[464] = inter_4[464];
    assign inter_5[465] = inter_4[465];
    assign inter_5[466] = inter_4[466];
    assign inter_5[467] = inter_4[467];
    assign inter_5[468] = inter_4[468];
    assign inter_5[469] = inter_4[469];
    assign inter_5[470] = inter_4[470];
    assign inter_5[471] = inter_4[471];
    assign inter_5[472] = inter_4[472];
    assign inter_5[473] = inter_4[473];
    assign inter_5[474] = inter_4[474];
    assign inter_5[475] = inter_4[475];
    assign inter_5[476] = inter_4[476];
    assign inter_5[477] = inter_4[477];
    assign inter_5[478] = inter_4[478];
    assign inter_5[479] = inter_4[479];
    assign inter_5[480] = inter_4[480]^inter_4[496];
    assign inter_5[481] = inter_4[481]^inter_4[497];
    assign inter_5[482] = inter_4[482]^inter_4[498];
    assign inter_5[483] = inter_4[483]^inter_4[499];
    assign inter_5[484] = inter_4[484]^inter_4[500];
    assign inter_5[485] = inter_4[485]^inter_4[501];
    assign inter_5[486] = inter_4[486]^inter_4[502];
    assign inter_5[487] = inter_4[487]^inter_4[503];
    assign inter_5[488] = inter_4[488]^inter_4[504];
    assign inter_5[489] = inter_4[489]^inter_4[505];
    assign inter_5[490] = inter_4[490]^inter_4[506];
    assign inter_5[491] = inter_4[491]^inter_4[507];
    assign inter_5[492] = inter_4[492]^inter_4[508];
    assign inter_5[493] = inter_4[493]^inter_4[509];
    assign inter_5[494] = inter_4[494]^inter_4[510];
    assign inter_5[495] = inter_4[495]^inter_4[511];
    assign inter_5[496] = inter_4[496];
    assign inter_5[497] = inter_4[497];
    assign inter_5[498] = inter_4[498];
    assign inter_5[499] = inter_4[499];
    assign inter_5[500] = inter_4[500];
    assign inter_5[501] = inter_4[501];
    assign inter_5[502] = inter_4[502];
    assign inter_5[503] = inter_4[503];
    assign inter_5[504] = inter_4[504];
    assign inter_5[505] = inter_4[505];
    assign inter_5[506] = inter_4[506];
    assign inter_5[507] = inter_4[507];
    assign inter_5[508] = inter_4[508];
    assign inter_5[509] = inter_4[509];
    assign inter_5[510] = inter_4[510];
    assign inter_5[511] = inter_4[511];
    assign inter_5[512] = inter_4[512]^inter_4[528];
    assign inter_5[513] = inter_4[513]^inter_4[529];
    assign inter_5[514] = inter_4[514]^inter_4[530];
    assign inter_5[515] = inter_4[515]^inter_4[531];
    assign inter_5[516] = inter_4[516]^inter_4[532];
    assign inter_5[517] = inter_4[517]^inter_4[533];
    assign inter_5[518] = inter_4[518]^inter_4[534];
    assign inter_5[519] = inter_4[519]^inter_4[535];
    assign inter_5[520] = inter_4[520]^inter_4[536];
    assign inter_5[521] = inter_4[521]^inter_4[537];
    assign inter_5[522] = inter_4[522]^inter_4[538];
    assign inter_5[523] = inter_4[523]^inter_4[539];
    assign inter_5[524] = inter_4[524]^inter_4[540];
    assign inter_5[525] = inter_4[525]^inter_4[541];
    assign inter_5[526] = inter_4[526]^inter_4[542];
    assign inter_5[527] = inter_4[527]^inter_4[543];
    assign inter_5[528] = inter_4[528];
    assign inter_5[529] = inter_4[529];
    assign inter_5[530] = inter_4[530];
    assign inter_5[531] = inter_4[531];
    assign inter_5[532] = inter_4[532];
    assign inter_5[533] = inter_4[533];
    assign inter_5[534] = inter_4[534];
    assign inter_5[535] = inter_4[535];
    assign inter_5[536] = inter_4[536];
    assign inter_5[537] = inter_4[537];
    assign inter_5[538] = inter_4[538];
    assign inter_5[539] = inter_4[539];
    assign inter_5[540] = inter_4[540];
    assign inter_5[541] = inter_4[541];
    assign inter_5[542] = inter_4[542];
    assign inter_5[543] = inter_4[543];
    assign inter_5[544] = inter_4[544]^inter_4[560];
    assign inter_5[545] = inter_4[545]^inter_4[561];
    assign inter_5[546] = inter_4[546]^inter_4[562];
    assign inter_5[547] = inter_4[547]^inter_4[563];
    assign inter_5[548] = inter_4[548]^inter_4[564];
    assign inter_5[549] = inter_4[549]^inter_4[565];
    assign inter_5[550] = inter_4[550]^inter_4[566];
    assign inter_5[551] = inter_4[551]^inter_4[567];
    assign inter_5[552] = inter_4[552]^inter_4[568];
    assign inter_5[553] = inter_4[553]^inter_4[569];
    assign inter_5[554] = inter_4[554]^inter_4[570];
    assign inter_5[555] = inter_4[555]^inter_4[571];
    assign inter_5[556] = inter_4[556]^inter_4[572];
    assign inter_5[557] = inter_4[557]^inter_4[573];
    assign inter_5[558] = inter_4[558]^inter_4[574];
    assign inter_5[559] = inter_4[559]^inter_4[575];
    assign inter_5[560] = inter_4[560];
    assign inter_5[561] = inter_4[561];
    assign inter_5[562] = inter_4[562];
    assign inter_5[563] = inter_4[563];
    assign inter_5[564] = inter_4[564];
    assign inter_5[565] = inter_4[565];
    assign inter_5[566] = inter_4[566];
    assign inter_5[567] = inter_4[567];
    assign inter_5[568] = inter_4[568];
    assign inter_5[569] = inter_4[569];
    assign inter_5[570] = inter_4[570];
    assign inter_5[571] = inter_4[571];
    assign inter_5[572] = inter_4[572];
    assign inter_5[573] = inter_4[573];
    assign inter_5[574] = inter_4[574];
    assign inter_5[575] = inter_4[575];
    assign inter_5[576] = inter_4[576]^inter_4[592];
    assign inter_5[577] = inter_4[577]^inter_4[593];
    assign inter_5[578] = inter_4[578]^inter_4[594];
    assign inter_5[579] = inter_4[579]^inter_4[595];
    assign inter_5[580] = inter_4[580]^inter_4[596];
    assign inter_5[581] = inter_4[581]^inter_4[597];
    assign inter_5[582] = inter_4[582]^inter_4[598];
    assign inter_5[583] = inter_4[583]^inter_4[599];
    assign inter_5[584] = inter_4[584]^inter_4[600];
    assign inter_5[585] = inter_4[585]^inter_4[601];
    assign inter_5[586] = inter_4[586]^inter_4[602];
    assign inter_5[587] = inter_4[587]^inter_4[603];
    assign inter_5[588] = inter_4[588]^inter_4[604];
    assign inter_5[589] = inter_4[589]^inter_4[605];
    assign inter_5[590] = inter_4[590]^inter_4[606];
    assign inter_5[591] = inter_4[591]^inter_4[607];
    assign inter_5[592] = inter_4[592];
    assign inter_5[593] = inter_4[593];
    assign inter_5[594] = inter_4[594];
    assign inter_5[595] = inter_4[595];
    assign inter_5[596] = inter_4[596];
    assign inter_5[597] = inter_4[597];
    assign inter_5[598] = inter_4[598];
    assign inter_5[599] = inter_4[599];
    assign inter_5[600] = inter_4[600];
    assign inter_5[601] = inter_4[601];
    assign inter_5[602] = inter_4[602];
    assign inter_5[603] = inter_4[603];
    assign inter_5[604] = inter_4[604];
    assign inter_5[605] = inter_4[605];
    assign inter_5[606] = inter_4[606];
    assign inter_5[607] = inter_4[607];
    assign inter_5[608] = inter_4[608]^inter_4[624];
    assign inter_5[609] = inter_4[609]^inter_4[625];
    assign inter_5[610] = inter_4[610]^inter_4[626];
    assign inter_5[611] = inter_4[611]^inter_4[627];
    assign inter_5[612] = inter_4[612]^inter_4[628];
    assign inter_5[613] = inter_4[613]^inter_4[629];
    assign inter_5[614] = inter_4[614]^inter_4[630];
    assign inter_5[615] = inter_4[615]^inter_4[631];
    assign inter_5[616] = inter_4[616]^inter_4[632];
    assign inter_5[617] = inter_4[617]^inter_4[633];
    assign inter_5[618] = inter_4[618]^inter_4[634];
    assign inter_5[619] = inter_4[619]^inter_4[635];
    assign inter_5[620] = inter_4[620]^inter_4[636];
    assign inter_5[621] = inter_4[621]^inter_4[637];
    assign inter_5[622] = inter_4[622]^inter_4[638];
    assign inter_5[623] = inter_4[623]^inter_4[639];
    assign inter_5[624] = inter_4[624];
    assign inter_5[625] = inter_4[625];
    assign inter_5[626] = inter_4[626];
    assign inter_5[627] = inter_4[627];
    assign inter_5[628] = inter_4[628];
    assign inter_5[629] = inter_4[629];
    assign inter_5[630] = inter_4[630];
    assign inter_5[631] = inter_4[631];
    assign inter_5[632] = inter_4[632];
    assign inter_5[633] = inter_4[633];
    assign inter_5[634] = inter_4[634];
    assign inter_5[635] = inter_4[635];
    assign inter_5[636] = inter_4[636];
    assign inter_5[637] = inter_4[637];
    assign inter_5[638] = inter_4[638];
    assign inter_5[639] = inter_4[639];
    assign inter_5[640] = inter_4[640]^inter_4[656];
    assign inter_5[641] = inter_4[641]^inter_4[657];
    assign inter_5[642] = inter_4[642]^inter_4[658];
    assign inter_5[643] = inter_4[643]^inter_4[659];
    assign inter_5[644] = inter_4[644]^inter_4[660];
    assign inter_5[645] = inter_4[645]^inter_4[661];
    assign inter_5[646] = inter_4[646]^inter_4[662];
    assign inter_5[647] = inter_4[647]^inter_4[663];
    assign inter_5[648] = inter_4[648]^inter_4[664];
    assign inter_5[649] = inter_4[649]^inter_4[665];
    assign inter_5[650] = inter_4[650]^inter_4[666];
    assign inter_5[651] = inter_4[651]^inter_4[667];
    assign inter_5[652] = inter_4[652]^inter_4[668];
    assign inter_5[653] = inter_4[653]^inter_4[669];
    assign inter_5[654] = inter_4[654]^inter_4[670];
    assign inter_5[655] = inter_4[655]^inter_4[671];
    assign inter_5[656] = inter_4[656];
    assign inter_5[657] = inter_4[657];
    assign inter_5[658] = inter_4[658];
    assign inter_5[659] = inter_4[659];
    assign inter_5[660] = inter_4[660];
    assign inter_5[661] = inter_4[661];
    assign inter_5[662] = inter_4[662];
    assign inter_5[663] = inter_4[663];
    assign inter_5[664] = inter_4[664];
    assign inter_5[665] = inter_4[665];
    assign inter_5[666] = inter_4[666];
    assign inter_5[667] = inter_4[667];
    assign inter_5[668] = inter_4[668];
    assign inter_5[669] = inter_4[669];
    assign inter_5[670] = inter_4[670];
    assign inter_5[671] = inter_4[671];
    assign inter_5[672] = inter_4[672]^inter_4[688];
    assign inter_5[673] = inter_4[673]^inter_4[689];
    assign inter_5[674] = inter_4[674]^inter_4[690];
    assign inter_5[675] = inter_4[675]^inter_4[691];
    assign inter_5[676] = inter_4[676]^inter_4[692];
    assign inter_5[677] = inter_4[677]^inter_4[693];
    assign inter_5[678] = inter_4[678]^inter_4[694];
    assign inter_5[679] = inter_4[679]^inter_4[695];
    assign inter_5[680] = inter_4[680]^inter_4[696];
    assign inter_5[681] = inter_4[681]^inter_4[697];
    assign inter_5[682] = inter_4[682]^inter_4[698];
    assign inter_5[683] = inter_4[683]^inter_4[699];
    assign inter_5[684] = inter_4[684]^inter_4[700];
    assign inter_5[685] = inter_4[685]^inter_4[701];
    assign inter_5[686] = inter_4[686]^inter_4[702];
    assign inter_5[687] = inter_4[687]^inter_4[703];
    assign inter_5[688] = inter_4[688];
    assign inter_5[689] = inter_4[689];
    assign inter_5[690] = inter_4[690];
    assign inter_5[691] = inter_4[691];
    assign inter_5[692] = inter_4[692];
    assign inter_5[693] = inter_4[693];
    assign inter_5[694] = inter_4[694];
    assign inter_5[695] = inter_4[695];
    assign inter_5[696] = inter_4[696];
    assign inter_5[697] = inter_4[697];
    assign inter_5[698] = inter_4[698];
    assign inter_5[699] = inter_4[699];
    assign inter_5[700] = inter_4[700];
    assign inter_5[701] = inter_4[701];
    assign inter_5[702] = inter_4[702];
    assign inter_5[703] = inter_4[703];
    assign inter_5[704] = inter_4[704]^inter_4[720];
    assign inter_5[705] = inter_4[705]^inter_4[721];
    assign inter_5[706] = inter_4[706]^inter_4[722];
    assign inter_5[707] = inter_4[707]^inter_4[723];
    assign inter_5[708] = inter_4[708]^inter_4[724];
    assign inter_5[709] = inter_4[709]^inter_4[725];
    assign inter_5[710] = inter_4[710]^inter_4[726];
    assign inter_5[711] = inter_4[711]^inter_4[727];
    assign inter_5[712] = inter_4[712]^inter_4[728];
    assign inter_5[713] = inter_4[713]^inter_4[729];
    assign inter_5[714] = inter_4[714]^inter_4[730];
    assign inter_5[715] = inter_4[715]^inter_4[731];
    assign inter_5[716] = inter_4[716]^inter_4[732];
    assign inter_5[717] = inter_4[717]^inter_4[733];
    assign inter_5[718] = inter_4[718]^inter_4[734];
    assign inter_5[719] = inter_4[719]^inter_4[735];
    assign inter_5[720] = inter_4[720];
    assign inter_5[721] = inter_4[721];
    assign inter_5[722] = inter_4[722];
    assign inter_5[723] = inter_4[723];
    assign inter_5[724] = inter_4[724];
    assign inter_5[725] = inter_4[725];
    assign inter_5[726] = inter_4[726];
    assign inter_5[727] = inter_4[727];
    assign inter_5[728] = inter_4[728];
    assign inter_5[729] = inter_4[729];
    assign inter_5[730] = inter_4[730];
    assign inter_5[731] = inter_4[731];
    assign inter_5[732] = inter_4[732];
    assign inter_5[733] = inter_4[733];
    assign inter_5[734] = inter_4[734];
    assign inter_5[735] = inter_4[735];
    assign inter_5[736] = inter_4[736]^inter_4[752];
    assign inter_5[737] = inter_4[737]^inter_4[753];
    assign inter_5[738] = inter_4[738]^inter_4[754];
    assign inter_5[739] = inter_4[739]^inter_4[755];
    assign inter_5[740] = inter_4[740]^inter_4[756];
    assign inter_5[741] = inter_4[741]^inter_4[757];
    assign inter_5[742] = inter_4[742]^inter_4[758];
    assign inter_5[743] = inter_4[743]^inter_4[759];
    assign inter_5[744] = inter_4[744]^inter_4[760];
    assign inter_5[745] = inter_4[745]^inter_4[761];
    assign inter_5[746] = inter_4[746]^inter_4[762];
    assign inter_5[747] = inter_4[747]^inter_4[763];
    assign inter_5[748] = inter_4[748]^inter_4[764];
    assign inter_5[749] = inter_4[749]^inter_4[765];
    assign inter_5[750] = inter_4[750]^inter_4[766];
    assign inter_5[751] = inter_4[751]^inter_4[767];
    assign inter_5[752] = inter_4[752];
    assign inter_5[753] = inter_4[753];
    assign inter_5[754] = inter_4[754];
    assign inter_5[755] = inter_4[755];
    assign inter_5[756] = inter_4[756];
    assign inter_5[757] = inter_4[757];
    assign inter_5[758] = inter_4[758];
    assign inter_5[759] = inter_4[759];
    assign inter_5[760] = inter_4[760];
    assign inter_5[761] = inter_4[761];
    assign inter_5[762] = inter_4[762];
    assign inter_5[763] = inter_4[763];
    assign inter_5[764] = inter_4[764];
    assign inter_5[765] = inter_4[765];
    assign inter_5[766] = inter_4[766];
    assign inter_5[767] = inter_4[767];
    assign inter_5[768] = inter_4[768]^inter_4[784];
    assign inter_5[769] = inter_4[769]^inter_4[785];
    assign inter_5[770] = inter_4[770]^inter_4[786];
    assign inter_5[771] = inter_4[771]^inter_4[787];
    assign inter_5[772] = inter_4[772]^inter_4[788];
    assign inter_5[773] = inter_4[773]^inter_4[789];
    assign inter_5[774] = inter_4[774]^inter_4[790];
    assign inter_5[775] = inter_4[775]^inter_4[791];
    assign inter_5[776] = inter_4[776]^inter_4[792];
    assign inter_5[777] = inter_4[777]^inter_4[793];
    assign inter_5[778] = inter_4[778]^inter_4[794];
    assign inter_5[779] = inter_4[779]^inter_4[795];
    assign inter_5[780] = inter_4[780]^inter_4[796];
    assign inter_5[781] = inter_4[781]^inter_4[797];
    assign inter_5[782] = inter_4[782]^inter_4[798];
    assign inter_5[783] = inter_4[783]^inter_4[799];
    assign inter_5[784] = inter_4[784];
    assign inter_5[785] = inter_4[785];
    assign inter_5[786] = inter_4[786];
    assign inter_5[787] = inter_4[787];
    assign inter_5[788] = inter_4[788];
    assign inter_5[789] = inter_4[789];
    assign inter_5[790] = inter_4[790];
    assign inter_5[791] = inter_4[791];
    assign inter_5[792] = inter_4[792];
    assign inter_5[793] = inter_4[793];
    assign inter_5[794] = inter_4[794];
    assign inter_5[795] = inter_4[795];
    assign inter_5[796] = inter_4[796];
    assign inter_5[797] = inter_4[797];
    assign inter_5[798] = inter_4[798];
    assign inter_5[799] = inter_4[799];
    assign inter_5[800] = inter_4[800]^inter_4[816];
    assign inter_5[801] = inter_4[801]^inter_4[817];
    assign inter_5[802] = inter_4[802]^inter_4[818];
    assign inter_5[803] = inter_4[803]^inter_4[819];
    assign inter_5[804] = inter_4[804]^inter_4[820];
    assign inter_5[805] = inter_4[805]^inter_4[821];
    assign inter_5[806] = inter_4[806]^inter_4[822];
    assign inter_5[807] = inter_4[807]^inter_4[823];
    assign inter_5[808] = inter_4[808]^inter_4[824];
    assign inter_5[809] = inter_4[809]^inter_4[825];
    assign inter_5[810] = inter_4[810]^inter_4[826];
    assign inter_5[811] = inter_4[811]^inter_4[827];
    assign inter_5[812] = inter_4[812]^inter_4[828];
    assign inter_5[813] = inter_4[813]^inter_4[829];
    assign inter_5[814] = inter_4[814]^inter_4[830];
    assign inter_5[815] = inter_4[815]^inter_4[831];
    assign inter_5[816] = inter_4[816];
    assign inter_5[817] = inter_4[817];
    assign inter_5[818] = inter_4[818];
    assign inter_5[819] = inter_4[819];
    assign inter_5[820] = inter_4[820];
    assign inter_5[821] = inter_4[821];
    assign inter_5[822] = inter_4[822];
    assign inter_5[823] = inter_4[823];
    assign inter_5[824] = inter_4[824];
    assign inter_5[825] = inter_4[825];
    assign inter_5[826] = inter_4[826];
    assign inter_5[827] = inter_4[827];
    assign inter_5[828] = inter_4[828];
    assign inter_5[829] = inter_4[829];
    assign inter_5[830] = inter_4[830];
    assign inter_5[831] = inter_4[831];
    assign inter_5[832] = inter_4[832]^inter_4[848];
    assign inter_5[833] = inter_4[833]^inter_4[849];
    assign inter_5[834] = inter_4[834]^inter_4[850];
    assign inter_5[835] = inter_4[835]^inter_4[851];
    assign inter_5[836] = inter_4[836]^inter_4[852];
    assign inter_5[837] = inter_4[837]^inter_4[853];
    assign inter_5[838] = inter_4[838]^inter_4[854];
    assign inter_5[839] = inter_4[839]^inter_4[855];
    assign inter_5[840] = inter_4[840]^inter_4[856];
    assign inter_5[841] = inter_4[841]^inter_4[857];
    assign inter_5[842] = inter_4[842]^inter_4[858];
    assign inter_5[843] = inter_4[843]^inter_4[859];
    assign inter_5[844] = inter_4[844]^inter_4[860];
    assign inter_5[845] = inter_4[845]^inter_4[861];
    assign inter_5[846] = inter_4[846]^inter_4[862];
    assign inter_5[847] = inter_4[847]^inter_4[863];
    assign inter_5[848] = inter_4[848];
    assign inter_5[849] = inter_4[849];
    assign inter_5[850] = inter_4[850];
    assign inter_5[851] = inter_4[851];
    assign inter_5[852] = inter_4[852];
    assign inter_5[853] = inter_4[853];
    assign inter_5[854] = inter_4[854];
    assign inter_5[855] = inter_4[855];
    assign inter_5[856] = inter_4[856];
    assign inter_5[857] = inter_4[857];
    assign inter_5[858] = inter_4[858];
    assign inter_5[859] = inter_4[859];
    assign inter_5[860] = inter_4[860];
    assign inter_5[861] = inter_4[861];
    assign inter_5[862] = inter_4[862];
    assign inter_5[863] = inter_4[863];
    assign inter_5[864] = inter_4[864]^inter_4[880];
    assign inter_5[865] = inter_4[865]^inter_4[881];
    assign inter_5[866] = inter_4[866]^inter_4[882];
    assign inter_5[867] = inter_4[867]^inter_4[883];
    assign inter_5[868] = inter_4[868]^inter_4[884];
    assign inter_5[869] = inter_4[869]^inter_4[885];
    assign inter_5[870] = inter_4[870]^inter_4[886];
    assign inter_5[871] = inter_4[871]^inter_4[887];
    assign inter_5[872] = inter_4[872]^inter_4[888];
    assign inter_5[873] = inter_4[873]^inter_4[889];
    assign inter_5[874] = inter_4[874]^inter_4[890];
    assign inter_5[875] = inter_4[875]^inter_4[891];
    assign inter_5[876] = inter_4[876]^inter_4[892];
    assign inter_5[877] = inter_4[877]^inter_4[893];
    assign inter_5[878] = inter_4[878]^inter_4[894];
    assign inter_5[879] = inter_4[879]^inter_4[895];
    assign inter_5[880] = inter_4[880];
    assign inter_5[881] = inter_4[881];
    assign inter_5[882] = inter_4[882];
    assign inter_5[883] = inter_4[883];
    assign inter_5[884] = inter_4[884];
    assign inter_5[885] = inter_4[885];
    assign inter_5[886] = inter_4[886];
    assign inter_5[887] = inter_4[887];
    assign inter_5[888] = inter_4[888];
    assign inter_5[889] = inter_4[889];
    assign inter_5[890] = inter_4[890];
    assign inter_5[891] = inter_4[891];
    assign inter_5[892] = inter_4[892];
    assign inter_5[893] = inter_4[893];
    assign inter_5[894] = inter_4[894];
    assign inter_5[895] = inter_4[895];
    assign inter_5[896] = inter_4[896]^inter_4[912];
    assign inter_5[897] = inter_4[897]^inter_4[913];
    assign inter_5[898] = inter_4[898]^inter_4[914];
    assign inter_5[899] = inter_4[899]^inter_4[915];
    assign inter_5[900] = inter_4[900]^inter_4[916];
    assign inter_5[901] = inter_4[901]^inter_4[917];
    assign inter_5[902] = inter_4[902]^inter_4[918];
    assign inter_5[903] = inter_4[903]^inter_4[919];
    assign inter_5[904] = inter_4[904]^inter_4[920];
    assign inter_5[905] = inter_4[905]^inter_4[921];
    assign inter_5[906] = inter_4[906]^inter_4[922];
    assign inter_5[907] = inter_4[907]^inter_4[923];
    assign inter_5[908] = inter_4[908]^inter_4[924];
    assign inter_5[909] = inter_4[909]^inter_4[925];
    assign inter_5[910] = inter_4[910]^inter_4[926];
    assign inter_5[911] = inter_4[911]^inter_4[927];
    assign inter_5[912] = inter_4[912];
    assign inter_5[913] = inter_4[913];
    assign inter_5[914] = inter_4[914];
    assign inter_5[915] = inter_4[915];
    assign inter_5[916] = inter_4[916];
    assign inter_5[917] = inter_4[917];
    assign inter_5[918] = inter_4[918];
    assign inter_5[919] = inter_4[919];
    assign inter_5[920] = inter_4[920];
    assign inter_5[921] = inter_4[921];
    assign inter_5[922] = inter_4[922];
    assign inter_5[923] = inter_4[923];
    assign inter_5[924] = inter_4[924];
    assign inter_5[925] = inter_4[925];
    assign inter_5[926] = inter_4[926];
    assign inter_5[927] = inter_4[927];
    assign inter_5[928] = inter_4[928]^inter_4[944];
    assign inter_5[929] = inter_4[929]^inter_4[945];
    assign inter_5[930] = inter_4[930]^inter_4[946];
    assign inter_5[931] = inter_4[931]^inter_4[947];
    assign inter_5[932] = inter_4[932]^inter_4[948];
    assign inter_5[933] = inter_4[933]^inter_4[949];
    assign inter_5[934] = inter_4[934]^inter_4[950];
    assign inter_5[935] = inter_4[935]^inter_4[951];
    assign inter_5[936] = inter_4[936]^inter_4[952];
    assign inter_5[937] = inter_4[937]^inter_4[953];
    assign inter_5[938] = inter_4[938]^inter_4[954];
    assign inter_5[939] = inter_4[939]^inter_4[955];
    assign inter_5[940] = inter_4[940]^inter_4[956];
    assign inter_5[941] = inter_4[941]^inter_4[957];
    assign inter_5[942] = inter_4[942]^inter_4[958];
    assign inter_5[943] = inter_4[943]^inter_4[959];
    assign inter_5[944] = inter_4[944];
    assign inter_5[945] = inter_4[945];
    assign inter_5[946] = inter_4[946];
    assign inter_5[947] = inter_4[947];
    assign inter_5[948] = inter_4[948];
    assign inter_5[949] = inter_4[949];
    assign inter_5[950] = inter_4[950];
    assign inter_5[951] = inter_4[951];
    assign inter_5[952] = inter_4[952];
    assign inter_5[953] = inter_4[953];
    assign inter_5[954] = inter_4[954];
    assign inter_5[955] = inter_4[955];
    assign inter_5[956] = inter_4[956];
    assign inter_5[957] = inter_4[957];
    assign inter_5[958] = inter_4[958];
    assign inter_5[959] = inter_4[959];
    assign inter_5[960] = inter_4[960]^inter_4[976];
    assign inter_5[961] = inter_4[961]^inter_4[977];
    assign inter_5[962] = inter_4[962]^inter_4[978];
    assign inter_5[963] = inter_4[963]^inter_4[979];
    assign inter_5[964] = inter_4[964]^inter_4[980];
    assign inter_5[965] = inter_4[965]^inter_4[981];
    assign inter_5[966] = inter_4[966]^inter_4[982];
    assign inter_5[967] = inter_4[967]^inter_4[983];
    assign inter_5[968] = inter_4[968]^inter_4[984];
    assign inter_5[969] = inter_4[969]^inter_4[985];
    assign inter_5[970] = inter_4[970]^inter_4[986];
    assign inter_5[971] = inter_4[971]^inter_4[987];
    assign inter_5[972] = inter_4[972]^inter_4[988];
    assign inter_5[973] = inter_4[973]^inter_4[989];
    assign inter_5[974] = inter_4[974]^inter_4[990];
    assign inter_5[975] = inter_4[975]^inter_4[991];
    assign inter_5[976] = inter_4[976];
    assign inter_5[977] = inter_4[977];
    assign inter_5[978] = inter_4[978];
    assign inter_5[979] = inter_4[979];
    assign inter_5[980] = inter_4[980];
    assign inter_5[981] = inter_4[981];
    assign inter_5[982] = inter_4[982];
    assign inter_5[983] = inter_4[983];
    assign inter_5[984] = inter_4[984];
    assign inter_5[985] = inter_4[985];
    assign inter_5[986] = inter_4[986];
    assign inter_5[987] = inter_4[987];
    assign inter_5[988] = inter_4[988];
    assign inter_5[989] = inter_4[989];
    assign inter_5[990] = inter_4[990];
    assign inter_5[991] = inter_4[991];
    assign inter_5[992] = inter_4[992]^inter_4[1008];
    assign inter_5[993] = inter_4[993]^inter_4[1009];
    assign inter_5[994] = inter_4[994]^inter_4[1010];
    assign inter_5[995] = inter_4[995]^inter_4[1011];
    assign inter_5[996] = inter_4[996]^inter_4[1012];
    assign inter_5[997] = inter_4[997]^inter_4[1013];
    assign inter_5[998] = inter_4[998]^inter_4[1014];
    assign inter_5[999] = inter_4[999]^inter_4[1015];
    assign inter_5[1000] = inter_4[1000]^inter_4[1016];
    assign inter_5[1001] = inter_4[1001]^inter_4[1017];
    assign inter_5[1002] = inter_4[1002]^inter_4[1018];
    assign inter_5[1003] = inter_4[1003]^inter_4[1019];
    assign inter_5[1004] = inter_4[1004]^inter_4[1020];
    assign inter_5[1005] = inter_4[1005]^inter_4[1021];
    assign inter_5[1006] = inter_4[1006]^inter_4[1022];
    assign inter_5[1007] = inter_4[1007]^inter_4[1023];
    assign inter_5[1008] = inter_4[1008];
    assign inter_5[1009] = inter_4[1009];
    assign inter_5[1010] = inter_4[1010];
    assign inter_5[1011] = inter_4[1011];
    assign inter_5[1012] = inter_4[1012];
    assign inter_5[1013] = inter_4[1013];
    assign inter_5[1014] = inter_4[1014];
    assign inter_5[1015] = inter_4[1015];
    assign inter_5[1016] = inter_4[1016];
    assign inter_5[1017] = inter_4[1017];
    assign inter_5[1018] = inter_4[1018];
    assign inter_5[1019] = inter_4[1019];
    assign inter_5[1020] = inter_4[1020];
    assign inter_5[1021] = inter_4[1021];
    assign inter_5[1022] = inter_4[1022];
    assign inter_5[1023] = inter_4[1023];
    /***************************/
    assign inter_6[0] = inter_5[0]^inter_5[32];
    assign inter_6[1] = inter_5[1]^inter_5[33];
    assign inter_6[2] = inter_5[2]^inter_5[34];
    assign inter_6[3] = inter_5[3]^inter_5[35];
    assign inter_6[4] = inter_5[4]^inter_5[36];
    assign inter_6[5] = inter_5[5]^inter_5[37];
    assign inter_6[6] = inter_5[6]^inter_5[38];
    assign inter_6[7] = inter_5[7]^inter_5[39];
    assign inter_6[8] = inter_5[8]^inter_5[40];
    assign inter_6[9] = inter_5[9]^inter_5[41];
    assign inter_6[10] = inter_5[10]^inter_5[42];
    assign inter_6[11] = inter_5[11]^inter_5[43];
    assign inter_6[12] = inter_5[12]^inter_5[44];
    assign inter_6[13] = inter_5[13]^inter_5[45];
    assign inter_6[14] = inter_5[14]^inter_5[46];
    assign inter_6[15] = inter_5[15]^inter_5[47];
    assign inter_6[16] = inter_5[16]^inter_5[48];
    assign inter_6[17] = inter_5[17]^inter_5[49];
    assign inter_6[18] = inter_5[18]^inter_5[50];
    assign inter_6[19] = inter_5[19]^inter_5[51];
    assign inter_6[20] = inter_5[20]^inter_5[52];
    assign inter_6[21] = inter_5[21]^inter_5[53];
    assign inter_6[22] = inter_5[22]^inter_5[54];
    assign inter_6[23] = inter_5[23]^inter_5[55];
    assign inter_6[24] = inter_5[24]^inter_5[56];
    assign inter_6[25] = inter_5[25]^inter_5[57];
    assign inter_6[26] = inter_5[26]^inter_5[58];
    assign inter_6[27] = inter_5[27]^inter_5[59];
    assign inter_6[28] = inter_5[28]^inter_5[60];
    assign inter_6[29] = inter_5[29]^inter_5[61];
    assign inter_6[30] = inter_5[30]^inter_5[62];
    assign inter_6[31] = inter_5[31]^inter_5[63];
    assign inter_6[32] = inter_5[32];
    assign inter_6[33] = inter_5[33];
    assign inter_6[34] = inter_5[34];
    assign inter_6[35] = inter_5[35];
    assign inter_6[36] = inter_5[36];
    assign inter_6[37] = inter_5[37];
    assign inter_6[38] = inter_5[38];
    assign inter_6[39] = inter_5[39];
    assign inter_6[40] = inter_5[40];
    assign inter_6[41] = inter_5[41];
    assign inter_6[42] = inter_5[42];
    assign inter_6[43] = inter_5[43];
    assign inter_6[44] = inter_5[44];
    assign inter_6[45] = inter_5[45];
    assign inter_6[46] = inter_5[46];
    assign inter_6[47] = inter_5[47];
    assign inter_6[48] = inter_5[48];
    assign inter_6[49] = inter_5[49];
    assign inter_6[50] = inter_5[50];
    assign inter_6[51] = inter_5[51];
    assign inter_6[52] = inter_5[52];
    assign inter_6[53] = inter_5[53];
    assign inter_6[54] = inter_5[54];
    assign inter_6[55] = inter_5[55];
    assign inter_6[56] = inter_5[56];
    assign inter_6[57] = inter_5[57];
    assign inter_6[58] = inter_5[58];
    assign inter_6[59] = inter_5[59];
    assign inter_6[60] = inter_5[60];
    assign inter_6[61] = inter_5[61];
    assign inter_6[62] = inter_5[62];
    assign inter_6[63] = inter_5[63];
    assign inter_6[64] = inter_5[64]^inter_5[96];
    assign inter_6[65] = inter_5[65]^inter_5[97];
    assign inter_6[66] = inter_5[66]^inter_5[98];
    assign inter_6[67] = inter_5[67]^inter_5[99];
    assign inter_6[68] = inter_5[68]^inter_5[100];
    assign inter_6[69] = inter_5[69]^inter_5[101];
    assign inter_6[70] = inter_5[70]^inter_5[102];
    assign inter_6[71] = inter_5[71]^inter_5[103];
    assign inter_6[72] = inter_5[72]^inter_5[104];
    assign inter_6[73] = inter_5[73]^inter_5[105];
    assign inter_6[74] = inter_5[74]^inter_5[106];
    assign inter_6[75] = inter_5[75]^inter_5[107];
    assign inter_6[76] = inter_5[76]^inter_5[108];
    assign inter_6[77] = inter_5[77]^inter_5[109];
    assign inter_6[78] = inter_5[78]^inter_5[110];
    assign inter_6[79] = inter_5[79]^inter_5[111];
    assign inter_6[80] = inter_5[80]^inter_5[112];
    assign inter_6[81] = inter_5[81]^inter_5[113];
    assign inter_6[82] = inter_5[82]^inter_5[114];
    assign inter_6[83] = inter_5[83]^inter_5[115];
    assign inter_6[84] = inter_5[84]^inter_5[116];
    assign inter_6[85] = inter_5[85]^inter_5[117];
    assign inter_6[86] = inter_5[86]^inter_5[118];
    assign inter_6[87] = inter_5[87]^inter_5[119];
    assign inter_6[88] = inter_5[88]^inter_5[120];
    assign inter_6[89] = inter_5[89]^inter_5[121];
    assign inter_6[90] = inter_5[90]^inter_5[122];
    assign inter_6[91] = inter_5[91]^inter_5[123];
    assign inter_6[92] = inter_5[92]^inter_5[124];
    assign inter_6[93] = inter_5[93]^inter_5[125];
    assign inter_6[94] = inter_5[94]^inter_5[126];
    assign inter_6[95] = inter_5[95]^inter_5[127];
    assign inter_6[96] = inter_5[96];
    assign inter_6[97] = inter_5[97];
    assign inter_6[98] = inter_5[98];
    assign inter_6[99] = inter_5[99];
    assign inter_6[100] = inter_5[100];
    assign inter_6[101] = inter_5[101];
    assign inter_6[102] = inter_5[102];
    assign inter_6[103] = inter_5[103];
    assign inter_6[104] = inter_5[104];
    assign inter_6[105] = inter_5[105];
    assign inter_6[106] = inter_5[106];
    assign inter_6[107] = inter_5[107];
    assign inter_6[108] = inter_5[108];
    assign inter_6[109] = inter_5[109];
    assign inter_6[110] = inter_5[110];
    assign inter_6[111] = inter_5[111];
    assign inter_6[112] = inter_5[112];
    assign inter_6[113] = inter_5[113];
    assign inter_6[114] = inter_5[114];
    assign inter_6[115] = inter_5[115];
    assign inter_6[116] = inter_5[116];
    assign inter_6[117] = inter_5[117];
    assign inter_6[118] = inter_5[118];
    assign inter_6[119] = inter_5[119];
    assign inter_6[120] = inter_5[120];
    assign inter_6[121] = inter_5[121];
    assign inter_6[122] = inter_5[122];
    assign inter_6[123] = inter_5[123];
    assign inter_6[124] = inter_5[124];
    assign inter_6[125] = inter_5[125];
    assign inter_6[126] = inter_5[126];
    assign inter_6[127] = inter_5[127];
    assign inter_6[128] = inter_5[128]^inter_5[160];
    assign inter_6[129] = inter_5[129]^inter_5[161];
    assign inter_6[130] = inter_5[130]^inter_5[162];
    assign inter_6[131] = inter_5[131]^inter_5[163];
    assign inter_6[132] = inter_5[132]^inter_5[164];
    assign inter_6[133] = inter_5[133]^inter_5[165];
    assign inter_6[134] = inter_5[134]^inter_5[166];
    assign inter_6[135] = inter_5[135]^inter_5[167];
    assign inter_6[136] = inter_5[136]^inter_5[168];
    assign inter_6[137] = inter_5[137]^inter_5[169];
    assign inter_6[138] = inter_5[138]^inter_5[170];
    assign inter_6[139] = inter_5[139]^inter_5[171];
    assign inter_6[140] = inter_5[140]^inter_5[172];
    assign inter_6[141] = inter_5[141]^inter_5[173];
    assign inter_6[142] = inter_5[142]^inter_5[174];
    assign inter_6[143] = inter_5[143]^inter_5[175];
    assign inter_6[144] = inter_5[144]^inter_5[176];
    assign inter_6[145] = inter_5[145]^inter_5[177];
    assign inter_6[146] = inter_5[146]^inter_5[178];
    assign inter_6[147] = inter_5[147]^inter_5[179];
    assign inter_6[148] = inter_5[148]^inter_5[180];
    assign inter_6[149] = inter_5[149]^inter_5[181];
    assign inter_6[150] = inter_5[150]^inter_5[182];
    assign inter_6[151] = inter_5[151]^inter_5[183];
    assign inter_6[152] = inter_5[152]^inter_5[184];
    assign inter_6[153] = inter_5[153]^inter_5[185];
    assign inter_6[154] = inter_5[154]^inter_5[186];
    assign inter_6[155] = inter_5[155]^inter_5[187];
    assign inter_6[156] = inter_5[156]^inter_5[188];
    assign inter_6[157] = inter_5[157]^inter_5[189];
    assign inter_6[158] = inter_5[158]^inter_5[190];
    assign inter_6[159] = inter_5[159]^inter_5[191];
    assign inter_6[160] = inter_5[160];
    assign inter_6[161] = inter_5[161];
    assign inter_6[162] = inter_5[162];
    assign inter_6[163] = inter_5[163];
    assign inter_6[164] = inter_5[164];
    assign inter_6[165] = inter_5[165];
    assign inter_6[166] = inter_5[166];
    assign inter_6[167] = inter_5[167];
    assign inter_6[168] = inter_5[168];
    assign inter_6[169] = inter_5[169];
    assign inter_6[170] = inter_5[170];
    assign inter_6[171] = inter_5[171];
    assign inter_6[172] = inter_5[172];
    assign inter_6[173] = inter_5[173];
    assign inter_6[174] = inter_5[174];
    assign inter_6[175] = inter_5[175];
    assign inter_6[176] = inter_5[176];
    assign inter_6[177] = inter_5[177];
    assign inter_6[178] = inter_5[178];
    assign inter_6[179] = inter_5[179];
    assign inter_6[180] = inter_5[180];
    assign inter_6[181] = inter_5[181];
    assign inter_6[182] = inter_5[182];
    assign inter_6[183] = inter_5[183];
    assign inter_6[184] = inter_5[184];
    assign inter_6[185] = inter_5[185];
    assign inter_6[186] = inter_5[186];
    assign inter_6[187] = inter_5[187];
    assign inter_6[188] = inter_5[188];
    assign inter_6[189] = inter_5[189];
    assign inter_6[190] = inter_5[190];
    assign inter_6[191] = inter_5[191];
    assign inter_6[192] = inter_5[192]^inter_5[224];
    assign inter_6[193] = inter_5[193]^inter_5[225];
    assign inter_6[194] = inter_5[194]^inter_5[226];
    assign inter_6[195] = inter_5[195]^inter_5[227];
    assign inter_6[196] = inter_5[196]^inter_5[228];
    assign inter_6[197] = inter_5[197]^inter_5[229];
    assign inter_6[198] = inter_5[198]^inter_5[230];
    assign inter_6[199] = inter_5[199]^inter_5[231];
    assign inter_6[200] = inter_5[200]^inter_5[232];
    assign inter_6[201] = inter_5[201]^inter_5[233];
    assign inter_6[202] = inter_5[202]^inter_5[234];
    assign inter_6[203] = inter_5[203]^inter_5[235];
    assign inter_6[204] = inter_5[204]^inter_5[236];
    assign inter_6[205] = inter_5[205]^inter_5[237];
    assign inter_6[206] = inter_5[206]^inter_5[238];
    assign inter_6[207] = inter_5[207]^inter_5[239];
    assign inter_6[208] = inter_5[208]^inter_5[240];
    assign inter_6[209] = inter_5[209]^inter_5[241];
    assign inter_6[210] = inter_5[210]^inter_5[242];
    assign inter_6[211] = inter_5[211]^inter_5[243];
    assign inter_6[212] = inter_5[212]^inter_5[244];
    assign inter_6[213] = inter_5[213]^inter_5[245];
    assign inter_6[214] = inter_5[214]^inter_5[246];
    assign inter_6[215] = inter_5[215]^inter_5[247];
    assign inter_6[216] = inter_5[216]^inter_5[248];
    assign inter_6[217] = inter_5[217]^inter_5[249];
    assign inter_6[218] = inter_5[218]^inter_5[250];
    assign inter_6[219] = inter_5[219]^inter_5[251];
    assign inter_6[220] = inter_5[220]^inter_5[252];
    assign inter_6[221] = inter_5[221]^inter_5[253];
    assign inter_6[222] = inter_5[222]^inter_5[254];
    assign inter_6[223] = inter_5[223]^inter_5[255];
    assign inter_6[224] = inter_5[224];
    assign inter_6[225] = inter_5[225];
    assign inter_6[226] = inter_5[226];
    assign inter_6[227] = inter_5[227];
    assign inter_6[228] = inter_5[228];
    assign inter_6[229] = inter_5[229];
    assign inter_6[230] = inter_5[230];
    assign inter_6[231] = inter_5[231];
    assign inter_6[232] = inter_5[232];
    assign inter_6[233] = inter_5[233];
    assign inter_6[234] = inter_5[234];
    assign inter_6[235] = inter_5[235];
    assign inter_6[236] = inter_5[236];
    assign inter_6[237] = inter_5[237];
    assign inter_6[238] = inter_5[238];
    assign inter_6[239] = inter_5[239];
    assign inter_6[240] = inter_5[240];
    assign inter_6[241] = inter_5[241];
    assign inter_6[242] = inter_5[242];
    assign inter_6[243] = inter_5[243];
    assign inter_6[244] = inter_5[244];
    assign inter_6[245] = inter_5[245];
    assign inter_6[246] = inter_5[246];
    assign inter_6[247] = inter_5[247];
    assign inter_6[248] = inter_5[248];
    assign inter_6[249] = inter_5[249];
    assign inter_6[250] = inter_5[250];
    assign inter_6[251] = inter_5[251];
    assign inter_6[252] = inter_5[252];
    assign inter_6[253] = inter_5[253];
    assign inter_6[254] = inter_5[254];
    assign inter_6[255] = inter_5[255];
    assign inter_6[256] = inter_5[256]^inter_5[288];
    assign inter_6[257] = inter_5[257]^inter_5[289];
    assign inter_6[258] = inter_5[258]^inter_5[290];
    assign inter_6[259] = inter_5[259]^inter_5[291];
    assign inter_6[260] = inter_5[260]^inter_5[292];
    assign inter_6[261] = inter_5[261]^inter_5[293];
    assign inter_6[262] = inter_5[262]^inter_5[294];
    assign inter_6[263] = inter_5[263]^inter_5[295];
    assign inter_6[264] = inter_5[264]^inter_5[296];
    assign inter_6[265] = inter_5[265]^inter_5[297];
    assign inter_6[266] = inter_5[266]^inter_5[298];
    assign inter_6[267] = inter_5[267]^inter_5[299];
    assign inter_6[268] = inter_5[268]^inter_5[300];
    assign inter_6[269] = inter_5[269]^inter_5[301];
    assign inter_6[270] = inter_5[270]^inter_5[302];
    assign inter_6[271] = inter_5[271]^inter_5[303];
    assign inter_6[272] = inter_5[272]^inter_5[304];
    assign inter_6[273] = inter_5[273]^inter_5[305];
    assign inter_6[274] = inter_5[274]^inter_5[306];
    assign inter_6[275] = inter_5[275]^inter_5[307];
    assign inter_6[276] = inter_5[276]^inter_5[308];
    assign inter_6[277] = inter_5[277]^inter_5[309];
    assign inter_6[278] = inter_5[278]^inter_5[310];
    assign inter_6[279] = inter_5[279]^inter_5[311];
    assign inter_6[280] = inter_5[280]^inter_5[312];
    assign inter_6[281] = inter_5[281]^inter_5[313];
    assign inter_6[282] = inter_5[282]^inter_5[314];
    assign inter_6[283] = inter_5[283]^inter_5[315];
    assign inter_6[284] = inter_5[284]^inter_5[316];
    assign inter_6[285] = inter_5[285]^inter_5[317];
    assign inter_6[286] = inter_5[286]^inter_5[318];
    assign inter_6[287] = inter_5[287]^inter_5[319];
    assign inter_6[288] = inter_5[288];
    assign inter_6[289] = inter_5[289];
    assign inter_6[290] = inter_5[290];
    assign inter_6[291] = inter_5[291];
    assign inter_6[292] = inter_5[292];
    assign inter_6[293] = inter_5[293];
    assign inter_6[294] = inter_5[294];
    assign inter_6[295] = inter_5[295];
    assign inter_6[296] = inter_5[296];
    assign inter_6[297] = inter_5[297];
    assign inter_6[298] = inter_5[298];
    assign inter_6[299] = inter_5[299];
    assign inter_6[300] = inter_5[300];
    assign inter_6[301] = inter_5[301];
    assign inter_6[302] = inter_5[302];
    assign inter_6[303] = inter_5[303];
    assign inter_6[304] = inter_5[304];
    assign inter_6[305] = inter_5[305];
    assign inter_6[306] = inter_5[306];
    assign inter_6[307] = inter_5[307];
    assign inter_6[308] = inter_5[308];
    assign inter_6[309] = inter_5[309];
    assign inter_6[310] = inter_5[310];
    assign inter_6[311] = inter_5[311];
    assign inter_6[312] = inter_5[312];
    assign inter_6[313] = inter_5[313];
    assign inter_6[314] = inter_5[314];
    assign inter_6[315] = inter_5[315];
    assign inter_6[316] = inter_5[316];
    assign inter_6[317] = inter_5[317];
    assign inter_6[318] = inter_5[318];
    assign inter_6[319] = inter_5[319];
    assign inter_6[320] = inter_5[320]^inter_5[352];
    assign inter_6[321] = inter_5[321]^inter_5[353];
    assign inter_6[322] = inter_5[322]^inter_5[354];
    assign inter_6[323] = inter_5[323]^inter_5[355];
    assign inter_6[324] = inter_5[324]^inter_5[356];
    assign inter_6[325] = inter_5[325]^inter_5[357];
    assign inter_6[326] = inter_5[326]^inter_5[358];
    assign inter_6[327] = inter_5[327]^inter_5[359];
    assign inter_6[328] = inter_5[328]^inter_5[360];
    assign inter_6[329] = inter_5[329]^inter_5[361];
    assign inter_6[330] = inter_5[330]^inter_5[362];
    assign inter_6[331] = inter_5[331]^inter_5[363];
    assign inter_6[332] = inter_5[332]^inter_5[364];
    assign inter_6[333] = inter_5[333]^inter_5[365];
    assign inter_6[334] = inter_5[334]^inter_5[366];
    assign inter_6[335] = inter_5[335]^inter_5[367];
    assign inter_6[336] = inter_5[336]^inter_5[368];
    assign inter_6[337] = inter_5[337]^inter_5[369];
    assign inter_6[338] = inter_5[338]^inter_5[370];
    assign inter_6[339] = inter_5[339]^inter_5[371];
    assign inter_6[340] = inter_5[340]^inter_5[372];
    assign inter_6[341] = inter_5[341]^inter_5[373];
    assign inter_6[342] = inter_5[342]^inter_5[374];
    assign inter_6[343] = inter_5[343]^inter_5[375];
    assign inter_6[344] = inter_5[344]^inter_5[376];
    assign inter_6[345] = inter_5[345]^inter_5[377];
    assign inter_6[346] = inter_5[346]^inter_5[378];
    assign inter_6[347] = inter_5[347]^inter_5[379];
    assign inter_6[348] = inter_5[348]^inter_5[380];
    assign inter_6[349] = inter_5[349]^inter_5[381];
    assign inter_6[350] = inter_5[350]^inter_5[382];
    assign inter_6[351] = inter_5[351]^inter_5[383];
    assign inter_6[352] = inter_5[352];
    assign inter_6[353] = inter_5[353];
    assign inter_6[354] = inter_5[354];
    assign inter_6[355] = inter_5[355];
    assign inter_6[356] = inter_5[356];
    assign inter_6[357] = inter_5[357];
    assign inter_6[358] = inter_5[358];
    assign inter_6[359] = inter_5[359];
    assign inter_6[360] = inter_5[360];
    assign inter_6[361] = inter_5[361];
    assign inter_6[362] = inter_5[362];
    assign inter_6[363] = inter_5[363];
    assign inter_6[364] = inter_5[364];
    assign inter_6[365] = inter_5[365];
    assign inter_6[366] = inter_5[366];
    assign inter_6[367] = inter_5[367];
    assign inter_6[368] = inter_5[368];
    assign inter_6[369] = inter_5[369];
    assign inter_6[370] = inter_5[370];
    assign inter_6[371] = inter_5[371];
    assign inter_6[372] = inter_5[372];
    assign inter_6[373] = inter_5[373];
    assign inter_6[374] = inter_5[374];
    assign inter_6[375] = inter_5[375];
    assign inter_6[376] = inter_5[376];
    assign inter_6[377] = inter_5[377];
    assign inter_6[378] = inter_5[378];
    assign inter_6[379] = inter_5[379];
    assign inter_6[380] = inter_5[380];
    assign inter_6[381] = inter_5[381];
    assign inter_6[382] = inter_5[382];
    assign inter_6[383] = inter_5[383];
    assign inter_6[384] = inter_5[384]^inter_5[416];
    assign inter_6[385] = inter_5[385]^inter_5[417];
    assign inter_6[386] = inter_5[386]^inter_5[418];
    assign inter_6[387] = inter_5[387]^inter_5[419];
    assign inter_6[388] = inter_5[388]^inter_5[420];
    assign inter_6[389] = inter_5[389]^inter_5[421];
    assign inter_6[390] = inter_5[390]^inter_5[422];
    assign inter_6[391] = inter_5[391]^inter_5[423];
    assign inter_6[392] = inter_5[392]^inter_5[424];
    assign inter_6[393] = inter_5[393]^inter_5[425];
    assign inter_6[394] = inter_5[394]^inter_5[426];
    assign inter_6[395] = inter_5[395]^inter_5[427];
    assign inter_6[396] = inter_5[396]^inter_5[428];
    assign inter_6[397] = inter_5[397]^inter_5[429];
    assign inter_6[398] = inter_5[398]^inter_5[430];
    assign inter_6[399] = inter_5[399]^inter_5[431];
    assign inter_6[400] = inter_5[400]^inter_5[432];
    assign inter_6[401] = inter_5[401]^inter_5[433];
    assign inter_6[402] = inter_5[402]^inter_5[434];
    assign inter_6[403] = inter_5[403]^inter_5[435];
    assign inter_6[404] = inter_5[404]^inter_5[436];
    assign inter_6[405] = inter_5[405]^inter_5[437];
    assign inter_6[406] = inter_5[406]^inter_5[438];
    assign inter_6[407] = inter_5[407]^inter_5[439];
    assign inter_6[408] = inter_5[408]^inter_5[440];
    assign inter_6[409] = inter_5[409]^inter_5[441];
    assign inter_6[410] = inter_5[410]^inter_5[442];
    assign inter_6[411] = inter_5[411]^inter_5[443];
    assign inter_6[412] = inter_5[412]^inter_5[444];
    assign inter_6[413] = inter_5[413]^inter_5[445];
    assign inter_6[414] = inter_5[414]^inter_5[446];
    assign inter_6[415] = inter_5[415]^inter_5[447];
    assign inter_6[416] = inter_5[416];
    assign inter_6[417] = inter_5[417];
    assign inter_6[418] = inter_5[418];
    assign inter_6[419] = inter_5[419];
    assign inter_6[420] = inter_5[420];
    assign inter_6[421] = inter_5[421];
    assign inter_6[422] = inter_5[422];
    assign inter_6[423] = inter_5[423];
    assign inter_6[424] = inter_5[424];
    assign inter_6[425] = inter_5[425];
    assign inter_6[426] = inter_5[426];
    assign inter_6[427] = inter_5[427];
    assign inter_6[428] = inter_5[428];
    assign inter_6[429] = inter_5[429];
    assign inter_6[430] = inter_5[430];
    assign inter_6[431] = inter_5[431];
    assign inter_6[432] = inter_5[432];
    assign inter_6[433] = inter_5[433];
    assign inter_6[434] = inter_5[434];
    assign inter_6[435] = inter_5[435];
    assign inter_6[436] = inter_5[436];
    assign inter_6[437] = inter_5[437];
    assign inter_6[438] = inter_5[438];
    assign inter_6[439] = inter_5[439];
    assign inter_6[440] = inter_5[440];
    assign inter_6[441] = inter_5[441];
    assign inter_6[442] = inter_5[442];
    assign inter_6[443] = inter_5[443];
    assign inter_6[444] = inter_5[444];
    assign inter_6[445] = inter_5[445];
    assign inter_6[446] = inter_5[446];
    assign inter_6[447] = inter_5[447];
    assign inter_6[448] = inter_5[448]^inter_5[480];
    assign inter_6[449] = inter_5[449]^inter_5[481];
    assign inter_6[450] = inter_5[450]^inter_5[482];
    assign inter_6[451] = inter_5[451]^inter_5[483];
    assign inter_6[452] = inter_5[452]^inter_5[484];
    assign inter_6[453] = inter_5[453]^inter_5[485];
    assign inter_6[454] = inter_5[454]^inter_5[486];
    assign inter_6[455] = inter_5[455]^inter_5[487];
    assign inter_6[456] = inter_5[456]^inter_5[488];
    assign inter_6[457] = inter_5[457]^inter_5[489];
    assign inter_6[458] = inter_5[458]^inter_5[490];
    assign inter_6[459] = inter_5[459]^inter_5[491];
    assign inter_6[460] = inter_5[460]^inter_5[492];
    assign inter_6[461] = inter_5[461]^inter_5[493];
    assign inter_6[462] = inter_5[462]^inter_5[494];
    assign inter_6[463] = inter_5[463]^inter_5[495];
    assign inter_6[464] = inter_5[464]^inter_5[496];
    assign inter_6[465] = inter_5[465]^inter_5[497];
    assign inter_6[466] = inter_5[466]^inter_5[498];
    assign inter_6[467] = inter_5[467]^inter_5[499];
    assign inter_6[468] = inter_5[468]^inter_5[500];
    assign inter_6[469] = inter_5[469]^inter_5[501];
    assign inter_6[470] = inter_5[470]^inter_5[502];
    assign inter_6[471] = inter_5[471]^inter_5[503];
    assign inter_6[472] = inter_5[472]^inter_5[504];
    assign inter_6[473] = inter_5[473]^inter_5[505];
    assign inter_6[474] = inter_5[474]^inter_5[506];
    assign inter_6[475] = inter_5[475]^inter_5[507];
    assign inter_6[476] = inter_5[476]^inter_5[508];
    assign inter_6[477] = inter_5[477]^inter_5[509];
    assign inter_6[478] = inter_5[478]^inter_5[510];
    assign inter_6[479] = inter_5[479]^inter_5[511];
    assign inter_6[480] = inter_5[480];
    assign inter_6[481] = inter_5[481];
    assign inter_6[482] = inter_5[482];
    assign inter_6[483] = inter_5[483];
    assign inter_6[484] = inter_5[484];
    assign inter_6[485] = inter_5[485];
    assign inter_6[486] = inter_5[486];
    assign inter_6[487] = inter_5[487];
    assign inter_6[488] = inter_5[488];
    assign inter_6[489] = inter_5[489];
    assign inter_6[490] = inter_5[490];
    assign inter_6[491] = inter_5[491];
    assign inter_6[492] = inter_5[492];
    assign inter_6[493] = inter_5[493];
    assign inter_6[494] = inter_5[494];
    assign inter_6[495] = inter_5[495];
    assign inter_6[496] = inter_5[496];
    assign inter_6[497] = inter_5[497];
    assign inter_6[498] = inter_5[498];
    assign inter_6[499] = inter_5[499];
    assign inter_6[500] = inter_5[500];
    assign inter_6[501] = inter_5[501];
    assign inter_6[502] = inter_5[502];
    assign inter_6[503] = inter_5[503];
    assign inter_6[504] = inter_5[504];
    assign inter_6[505] = inter_5[505];
    assign inter_6[506] = inter_5[506];
    assign inter_6[507] = inter_5[507];
    assign inter_6[508] = inter_5[508];
    assign inter_6[509] = inter_5[509];
    assign inter_6[510] = inter_5[510];
    assign inter_6[511] = inter_5[511];
    assign inter_6[512] = inter_5[512]^inter_5[544];
    assign inter_6[513] = inter_5[513]^inter_5[545];
    assign inter_6[514] = inter_5[514]^inter_5[546];
    assign inter_6[515] = inter_5[515]^inter_5[547];
    assign inter_6[516] = inter_5[516]^inter_5[548];
    assign inter_6[517] = inter_5[517]^inter_5[549];
    assign inter_6[518] = inter_5[518]^inter_5[550];
    assign inter_6[519] = inter_5[519]^inter_5[551];
    assign inter_6[520] = inter_5[520]^inter_5[552];
    assign inter_6[521] = inter_5[521]^inter_5[553];
    assign inter_6[522] = inter_5[522]^inter_5[554];
    assign inter_6[523] = inter_5[523]^inter_5[555];
    assign inter_6[524] = inter_5[524]^inter_5[556];
    assign inter_6[525] = inter_5[525]^inter_5[557];
    assign inter_6[526] = inter_5[526]^inter_5[558];
    assign inter_6[527] = inter_5[527]^inter_5[559];
    assign inter_6[528] = inter_5[528]^inter_5[560];
    assign inter_6[529] = inter_5[529]^inter_5[561];
    assign inter_6[530] = inter_5[530]^inter_5[562];
    assign inter_6[531] = inter_5[531]^inter_5[563];
    assign inter_6[532] = inter_5[532]^inter_5[564];
    assign inter_6[533] = inter_5[533]^inter_5[565];
    assign inter_6[534] = inter_5[534]^inter_5[566];
    assign inter_6[535] = inter_5[535]^inter_5[567];
    assign inter_6[536] = inter_5[536]^inter_5[568];
    assign inter_6[537] = inter_5[537]^inter_5[569];
    assign inter_6[538] = inter_5[538]^inter_5[570];
    assign inter_6[539] = inter_5[539]^inter_5[571];
    assign inter_6[540] = inter_5[540]^inter_5[572];
    assign inter_6[541] = inter_5[541]^inter_5[573];
    assign inter_6[542] = inter_5[542]^inter_5[574];
    assign inter_6[543] = inter_5[543]^inter_5[575];
    assign inter_6[544] = inter_5[544];
    assign inter_6[545] = inter_5[545];
    assign inter_6[546] = inter_5[546];
    assign inter_6[547] = inter_5[547];
    assign inter_6[548] = inter_5[548];
    assign inter_6[549] = inter_5[549];
    assign inter_6[550] = inter_5[550];
    assign inter_6[551] = inter_5[551];
    assign inter_6[552] = inter_5[552];
    assign inter_6[553] = inter_5[553];
    assign inter_6[554] = inter_5[554];
    assign inter_6[555] = inter_5[555];
    assign inter_6[556] = inter_5[556];
    assign inter_6[557] = inter_5[557];
    assign inter_6[558] = inter_5[558];
    assign inter_6[559] = inter_5[559];
    assign inter_6[560] = inter_5[560];
    assign inter_6[561] = inter_5[561];
    assign inter_6[562] = inter_5[562];
    assign inter_6[563] = inter_5[563];
    assign inter_6[564] = inter_5[564];
    assign inter_6[565] = inter_5[565];
    assign inter_6[566] = inter_5[566];
    assign inter_6[567] = inter_5[567];
    assign inter_6[568] = inter_5[568];
    assign inter_6[569] = inter_5[569];
    assign inter_6[570] = inter_5[570];
    assign inter_6[571] = inter_5[571];
    assign inter_6[572] = inter_5[572];
    assign inter_6[573] = inter_5[573];
    assign inter_6[574] = inter_5[574];
    assign inter_6[575] = inter_5[575];
    assign inter_6[576] = inter_5[576]^inter_5[608];
    assign inter_6[577] = inter_5[577]^inter_5[609];
    assign inter_6[578] = inter_5[578]^inter_5[610];
    assign inter_6[579] = inter_5[579]^inter_5[611];
    assign inter_6[580] = inter_5[580]^inter_5[612];
    assign inter_6[581] = inter_5[581]^inter_5[613];
    assign inter_6[582] = inter_5[582]^inter_5[614];
    assign inter_6[583] = inter_5[583]^inter_5[615];
    assign inter_6[584] = inter_5[584]^inter_5[616];
    assign inter_6[585] = inter_5[585]^inter_5[617];
    assign inter_6[586] = inter_5[586]^inter_5[618];
    assign inter_6[587] = inter_5[587]^inter_5[619];
    assign inter_6[588] = inter_5[588]^inter_5[620];
    assign inter_6[589] = inter_5[589]^inter_5[621];
    assign inter_6[590] = inter_5[590]^inter_5[622];
    assign inter_6[591] = inter_5[591]^inter_5[623];
    assign inter_6[592] = inter_5[592]^inter_5[624];
    assign inter_6[593] = inter_5[593]^inter_5[625];
    assign inter_6[594] = inter_5[594]^inter_5[626];
    assign inter_6[595] = inter_5[595]^inter_5[627];
    assign inter_6[596] = inter_5[596]^inter_5[628];
    assign inter_6[597] = inter_5[597]^inter_5[629];
    assign inter_6[598] = inter_5[598]^inter_5[630];
    assign inter_6[599] = inter_5[599]^inter_5[631];
    assign inter_6[600] = inter_5[600]^inter_5[632];
    assign inter_6[601] = inter_5[601]^inter_5[633];
    assign inter_6[602] = inter_5[602]^inter_5[634];
    assign inter_6[603] = inter_5[603]^inter_5[635];
    assign inter_6[604] = inter_5[604]^inter_5[636];
    assign inter_6[605] = inter_5[605]^inter_5[637];
    assign inter_6[606] = inter_5[606]^inter_5[638];
    assign inter_6[607] = inter_5[607]^inter_5[639];
    assign inter_6[608] = inter_5[608];
    assign inter_6[609] = inter_5[609];
    assign inter_6[610] = inter_5[610];
    assign inter_6[611] = inter_5[611];
    assign inter_6[612] = inter_5[612];
    assign inter_6[613] = inter_5[613];
    assign inter_6[614] = inter_5[614];
    assign inter_6[615] = inter_5[615];
    assign inter_6[616] = inter_5[616];
    assign inter_6[617] = inter_5[617];
    assign inter_6[618] = inter_5[618];
    assign inter_6[619] = inter_5[619];
    assign inter_6[620] = inter_5[620];
    assign inter_6[621] = inter_5[621];
    assign inter_6[622] = inter_5[622];
    assign inter_6[623] = inter_5[623];
    assign inter_6[624] = inter_5[624];
    assign inter_6[625] = inter_5[625];
    assign inter_6[626] = inter_5[626];
    assign inter_6[627] = inter_5[627];
    assign inter_6[628] = inter_5[628];
    assign inter_6[629] = inter_5[629];
    assign inter_6[630] = inter_5[630];
    assign inter_6[631] = inter_5[631];
    assign inter_6[632] = inter_5[632];
    assign inter_6[633] = inter_5[633];
    assign inter_6[634] = inter_5[634];
    assign inter_6[635] = inter_5[635];
    assign inter_6[636] = inter_5[636];
    assign inter_6[637] = inter_5[637];
    assign inter_6[638] = inter_5[638];
    assign inter_6[639] = inter_5[639];
    assign inter_6[640] = inter_5[640]^inter_5[672];
    assign inter_6[641] = inter_5[641]^inter_5[673];
    assign inter_6[642] = inter_5[642]^inter_5[674];
    assign inter_6[643] = inter_5[643]^inter_5[675];
    assign inter_6[644] = inter_5[644]^inter_5[676];
    assign inter_6[645] = inter_5[645]^inter_5[677];
    assign inter_6[646] = inter_5[646]^inter_5[678];
    assign inter_6[647] = inter_5[647]^inter_5[679];
    assign inter_6[648] = inter_5[648]^inter_5[680];
    assign inter_6[649] = inter_5[649]^inter_5[681];
    assign inter_6[650] = inter_5[650]^inter_5[682];
    assign inter_6[651] = inter_5[651]^inter_5[683];
    assign inter_6[652] = inter_5[652]^inter_5[684];
    assign inter_6[653] = inter_5[653]^inter_5[685];
    assign inter_6[654] = inter_5[654]^inter_5[686];
    assign inter_6[655] = inter_5[655]^inter_5[687];
    assign inter_6[656] = inter_5[656]^inter_5[688];
    assign inter_6[657] = inter_5[657]^inter_5[689];
    assign inter_6[658] = inter_5[658]^inter_5[690];
    assign inter_6[659] = inter_5[659]^inter_5[691];
    assign inter_6[660] = inter_5[660]^inter_5[692];
    assign inter_6[661] = inter_5[661]^inter_5[693];
    assign inter_6[662] = inter_5[662]^inter_5[694];
    assign inter_6[663] = inter_5[663]^inter_5[695];
    assign inter_6[664] = inter_5[664]^inter_5[696];
    assign inter_6[665] = inter_5[665]^inter_5[697];
    assign inter_6[666] = inter_5[666]^inter_5[698];
    assign inter_6[667] = inter_5[667]^inter_5[699];
    assign inter_6[668] = inter_5[668]^inter_5[700];
    assign inter_6[669] = inter_5[669]^inter_5[701];
    assign inter_6[670] = inter_5[670]^inter_5[702];
    assign inter_6[671] = inter_5[671]^inter_5[703];
    assign inter_6[672] = inter_5[672];
    assign inter_6[673] = inter_5[673];
    assign inter_6[674] = inter_5[674];
    assign inter_6[675] = inter_5[675];
    assign inter_6[676] = inter_5[676];
    assign inter_6[677] = inter_5[677];
    assign inter_6[678] = inter_5[678];
    assign inter_6[679] = inter_5[679];
    assign inter_6[680] = inter_5[680];
    assign inter_6[681] = inter_5[681];
    assign inter_6[682] = inter_5[682];
    assign inter_6[683] = inter_5[683];
    assign inter_6[684] = inter_5[684];
    assign inter_6[685] = inter_5[685];
    assign inter_6[686] = inter_5[686];
    assign inter_6[687] = inter_5[687];
    assign inter_6[688] = inter_5[688];
    assign inter_6[689] = inter_5[689];
    assign inter_6[690] = inter_5[690];
    assign inter_6[691] = inter_5[691];
    assign inter_6[692] = inter_5[692];
    assign inter_6[693] = inter_5[693];
    assign inter_6[694] = inter_5[694];
    assign inter_6[695] = inter_5[695];
    assign inter_6[696] = inter_5[696];
    assign inter_6[697] = inter_5[697];
    assign inter_6[698] = inter_5[698];
    assign inter_6[699] = inter_5[699];
    assign inter_6[700] = inter_5[700];
    assign inter_6[701] = inter_5[701];
    assign inter_6[702] = inter_5[702];
    assign inter_6[703] = inter_5[703];
    assign inter_6[704] = inter_5[704]^inter_5[736];
    assign inter_6[705] = inter_5[705]^inter_5[737];
    assign inter_6[706] = inter_5[706]^inter_5[738];
    assign inter_6[707] = inter_5[707]^inter_5[739];
    assign inter_6[708] = inter_5[708]^inter_5[740];
    assign inter_6[709] = inter_5[709]^inter_5[741];
    assign inter_6[710] = inter_5[710]^inter_5[742];
    assign inter_6[711] = inter_5[711]^inter_5[743];
    assign inter_6[712] = inter_5[712]^inter_5[744];
    assign inter_6[713] = inter_5[713]^inter_5[745];
    assign inter_6[714] = inter_5[714]^inter_5[746];
    assign inter_6[715] = inter_5[715]^inter_5[747];
    assign inter_6[716] = inter_5[716]^inter_5[748];
    assign inter_6[717] = inter_5[717]^inter_5[749];
    assign inter_6[718] = inter_5[718]^inter_5[750];
    assign inter_6[719] = inter_5[719]^inter_5[751];
    assign inter_6[720] = inter_5[720]^inter_5[752];
    assign inter_6[721] = inter_5[721]^inter_5[753];
    assign inter_6[722] = inter_5[722]^inter_5[754];
    assign inter_6[723] = inter_5[723]^inter_5[755];
    assign inter_6[724] = inter_5[724]^inter_5[756];
    assign inter_6[725] = inter_5[725]^inter_5[757];
    assign inter_6[726] = inter_5[726]^inter_5[758];
    assign inter_6[727] = inter_5[727]^inter_5[759];
    assign inter_6[728] = inter_5[728]^inter_5[760];
    assign inter_6[729] = inter_5[729]^inter_5[761];
    assign inter_6[730] = inter_5[730]^inter_5[762];
    assign inter_6[731] = inter_5[731]^inter_5[763];
    assign inter_6[732] = inter_5[732]^inter_5[764];
    assign inter_6[733] = inter_5[733]^inter_5[765];
    assign inter_6[734] = inter_5[734]^inter_5[766];
    assign inter_6[735] = inter_5[735]^inter_5[767];
    assign inter_6[736] = inter_5[736];
    assign inter_6[737] = inter_5[737];
    assign inter_6[738] = inter_5[738];
    assign inter_6[739] = inter_5[739];
    assign inter_6[740] = inter_5[740];
    assign inter_6[741] = inter_5[741];
    assign inter_6[742] = inter_5[742];
    assign inter_6[743] = inter_5[743];
    assign inter_6[744] = inter_5[744];
    assign inter_6[745] = inter_5[745];
    assign inter_6[746] = inter_5[746];
    assign inter_6[747] = inter_5[747];
    assign inter_6[748] = inter_5[748];
    assign inter_6[749] = inter_5[749];
    assign inter_6[750] = inter_5[750];
    assign inter_6[751] = inter_5[751];
    assign inter_6[752] = inter_5[752];
    assign inter_6[753] = inter_5[753];
    assign inter_6[754] = inter_5[754];
    assign inter_6[755] = inter_5[755];
    assign inter_6[756] = inter_5[756];
    assign inter_6[757] = inter_5[757];
    assign inter_6[758] = inter_5[758];
    assign inter_6[759] = inter_5[759];
    assign inter_6[760] = inter_5[760];
    assign inter_6[761] = inter_5[761];
    assign inter_6[762] = inter_5[762];
    assign inter_6[763] = inter_5[763];
    assign inter_6[764] = inter_5[764];
    assign inter_6[765] = inter_5[765];
    assign inter_6[766] = inter_5[766];
    assign inter_6[767] = inter_5[767];
    assign inter_6[768] = inter_5[768]^inter_5[800];
    assign inter_6[769] = inter_5[769]^inter_5[801];
    assign inter_6[770] = inter_5[770]^inter_5[802];
    assign inter_6[771] = inter_5[771]^inter_5[803];
    assign inter_6[772] = inter_5[772]^inter_5[804];
    assign inter_6[773] = inter_5[773]^inter_5[805];
    assign inter_6[774] = inter_5[774]^inter_5[806];
    assign inter_6[775] = inter_5[775]^inter_5[807];
    assign inter_6[776] = inter_5[776]^inter_5[808];
    assign inter_6[777] = inter_5[777]^inter_5[809];
    assign inter_6[778] = inter_5[778]^inter_5[810];
    assign inter_6[779] = inter_5[779]^inter_5[811];
    assign inter_6[780] = inter_5[780]^inter_5[812];
    assign inter_6[781] = inter_5[781]^inter_5[813];
    assign inter_6[782] = inter_5[782]^inter_5[814];
    assign inter_6[783] = inter_5[783]^inter_5[815];
    assign inter_6[784] = inter_5[784]^inter_5[816];
    assign inter_6[785] = inter_5[785]^inter_5[817];
    assign inter_6[786] = inter_5[786]^inter_5[818];
    assign inter_6[787] = inter_5[787]^inter_5[819];
    assign inter_6[788] = inter_5[788]^inter_5[820];
    assign inter_6[789] = inter_5[789]^inter_5[821];
    assign inter_6[790] = inter_5[790]^inter_5[822];
    assign inter_6[791] = inter_5[791]^inter_5[823];
    assign inter_6[792] = inter_5[792]^inter_5[824];
    assign inter_6[793] = inter_5[793]^inter_5[825];
    assign inter_6[794] = inter_5[794]^inter_5[826];
    assign inter_6[795] = inter_5[795]^inter_5[827];
    assign inter_6[796] = inter_5[796]^inter_5[828];
    assign inter_6[797] = inter_5[797]^inter_5[829];
    assign inter_6[798] = inter_5[798]^inter_5[830];
    assign inter_6[799] = inter_5[799]^inter_5[831];
    assign inter_6[800] = inter_5[800];
    assign inter_6[801] = inter_5[801];
    assign inter_6[802] = inter_5[802];
    assign inter_6[803] = inter_5[803];
    assign inter_6[804] = inter_5[804];
    assign inter_6[805] = inter_5[805];
    assign inter_6[806] = inter_5[806];
    assign inter_6[807] = inter_5[807];
    assign inter_6[808] = inter_5[808];
    assign inter_6[809] = inter_5[809];
    assign inter_6[810] = inter_5[810];
    assign inter_6[811] = inter_5[811];
    assign inter_6[812] = inter_5[812];
    assign inter_6[813] = inter_5[813];
    assign inter_6[814] = inter_5[814];
    assign inter_6[815] = inter_5[815];
    assign inter_6[816] = inter_5[816];
    assign inter_6[817] = inter_5[817];
    assign inter_6[818] = inter_5[818];
    assign inter_6[819] = inter_5[819];
    assign inter_6[820] = inter_5[820];
    assign inter_6[821] = inter_5[821];
    assign inter_6[822] = inter_5[822];
    assign inter_6[823] = inter_5[823];
    assign inter_6[824] = inter_5[824];
    assign inter_6[825] = inter_5[825];
    assign inter_6[826] = inter_5[826];
    assign inter_6[827] = inter_5[827];
    assign inter_6[828] = inter_5[828];
    assign inter_6[829] = inter_5[829];
    assign inter_6[830] = inter_5[830];
    assign inter_6[831] = inter_5[831];
    assign inter_6[832] = inter_5[832]^inter_5[864];
    assign inter_6[833] = inter_5[833]^inter_5[865];
    assign inter_6[834] = inter_5[834]^inter_5[866];
    assign inter_6[835] = inter_5[835]^inter_5[867];
    assign inter_6[836] = inter_5[836]^inter_5[868];
    assign inter_6[837] = inter_5[837]^inter_5[869];
    assign inter_6[838] = inter_5[838]^inter_5[870];
    assign inter_6[839] = inter_5[839]^inter_5[871];
    assign inter_6[840] = inter_5[840]^inter_5[872];
    assign inter_6[841] = inter_5[841]^inter_5[873];
    assign inter_6[842] = inter_5[842]^inter_5[874];
    assign inter_6[843] = inter_5[843]^inter_5[875];
    assign inter_6[844] = inter_5[844]^inter_5[876];
    assign inter_6[845] = inter_5[845]^inter_5[877];
    assign inter_6[846] = inter_5[846]^inter_5[878];
    assign inter_6[847] = inter_5[847]^inter_5[879];
    assign inter_6[848] = inter_5[848]^inter_5[880];
    assign inter_6[849] = inter_5[849]^inter_5[881];
    assign inter_6[850] = inter_5[850]^inter_5[882];
    assign inter_6[851] = inter_5[851]^inter_5[883];
    assign inter_6[852] = inter_5[852]^inter_5[884];
    assign inter_6[853] = inter_5[853]^inter_5[885];
    assign inter_6[854] = inter_5[854]^inter_5[886];
    assign inter_6[855] = inter_5[855]^inter_5[887];
    assign inter_6[856] = inter_5[856]^inter_5[888];
    assign inter_6[857] = inter_5[857]^inter_5[889];
    assign inter_6[858] = inter_5[858]^inter_5[890];
    assign inter_6[859] = inter_5[859]^inter_5[891];
    assign inter_6[860] = inter_5[860]^inter_5[892];
    assign inter_6[861] = inter_5[861]^inter_5[893];
    assign inter_6[862] = inter_5[862]^inter_5[894];
    assign inter_6[863] = inter_5[863]^inter_5[895];
    assign inter_6[864] = inter_5[864];
    assign inter_6[865] = inter_5[865];
    assign inter_6[866] = inter_5[866];
    assign inter_6[867] = inter_5[867];
    assign inter_6[868] = inter_5[868];
    assign inter_6[869] = inter_5[869];
    assign inter_6[870] = inter_5[870];
    assign inter_6[871] = inter_5[871];
    assign inter_6[872] = inter_5[872];
    assign inter_6[873] = inter_5[873];
    assign inter_6[874] = inter_5[874];
    assign inter_6[875] = inter_5[875];
    assign inter_6[876] = inter_5[876];
    assign inter_6[877] = inter_5[877];
    assign inter_6[878] = inter_5[878];
    assign inter_6[879] = inter_5[879];
    assign inter_6[880] = inter_5[880];
    assign inter_6[881] = inter_5[881];
    assign inter_6[882] = inter_5[882];
    assign inter_6[883] = inter_5[883];
    assign inter_6[884] = inter_5[884];
    assign inter_6[885] = inter_5[885];
    assign inter_6[886] = inter_5[886];
    assign inter_6[887] = inter_5[887];
    assign inter_6[888] = inter_5[888];
    assign inter_6[889] = inter_5[889];
    assign inter_6[890] = inter_5[890];
    assign inter_6[891] = inter_5[891];
    assign inter_6[892] = inter_5[892];
    assign inter_6[893] = inter_5[893];
    assign inter_6[894] = inter_5[894];
    assign inter_6[895] = inter_5[895];
    assign inter_6[896] = inter_5[896]^inter_5[928];
    assign inter_6[897] = inter_5[897]^inter_5[929];
    assign inter_6[898] = inter_5[898]^inter_5[930];
    assign inter_6[899] = inter_5[899]^inter_5[931];
    assign inter_6[900] = inter_5[900]^inter_5[932];
    assign inter_6[901] = inter_5[901]^inter_5[933];
    assign inter_6[902] = inter_5[902]^inter_5[934];
    assign inter_6[903] = inter_5[903]^inter_5[935];
    assign inter_6[904] = inter_5[904]^inter_5[936];
    assign inter_6[905] = inter_5[905]^inter_5[937];
    assign inter_6[906] = inter_5[906]^inter_5[938];
    assign inter_6[907] = inter_5[907]^inter_5[939];
    assign inter_6[908] = inter_5[908]^inter_5[940];
    assign inter_6[909] = inter_5[909]^inter_5[941];
    assign inter_6[910] = inter_5[910]^inter_5[942];
    assign inter_6[911] = inter_5[911]^inter_5[943];
    assign inter_6[912] = inter_5[912]^inter_5[944];
    assign inter_6[913] = inter_5[913]^inter_5[945];
    assign inter_6[914] = inter_5[914]^inter_5[946];
    assign inter_6[915] = inter_5[915]^inter_5[947];
    assign inter_6[916] = inter_5[916]^inter_5[948];
    assign inter_6[917] = inter_5[917]^inter_5[949];
    assign inter_6[918] = inter_5[918]^inter_5[950];
    assign inter_6[919] = inter_5[919]^inter_5[951];
    assign inter_6[920] = inter_5[920]^inter_5[952];
    assign inter_6[921] = inter_5[921]^inter_5[953];
    assign inter_6[922] = inter_5[922]^inter_5[954];
    assign inter_6[923] = inter_5[923]^inter_5[955];
    assign inter_6[924] = inter_5[924]^inter_5[956];
    assign inter_6[925] = inter_5[925]^inter_5[957];
    assign inter_6[926] = inter_5[926]^inter_5[958];
    assign inter_6[927] = inter_5[927]^inter_5[959];
    assign inter_6[928] = inter_5[928];
    assign inter_6[929] = inter_5[929];
    assign inter_6[930] = inter_5[930];
    assign inter_6[931] = inter_5[931];
    assign inter_6[932] = inter_5[932];
    assign inter_6[933] = inter_5[933];
    assign inter_6[934] = inter_5[934];
    assign inter_6[935] = inter_5[935];
    assign inter_6[936] = inter_5[936];
    assign inter_6[937] = inter_5[937];
    assign inter_6[938] = inter_5[938];
    assign inter_6[939] = inter_5[939];
    assign inter_6[940] = inter_5[940];
    assign inter_6[941] = inter_5[941];
    assign inter_6[942] = inter_5[942];
    assign inter_6[943] = inter_5[943];
    assign inter_6[944] = inter_5[944];
    assign inter_6[945] = inter_5[945];
    assign inter_6[946] = inter_5[946];
    assign inter_6[947] = inter_5[947];
    assign inter_6[948] = inter_5[948];
    assign inter_6[949] = inter_5[949];
    assign inter_6[950] = inter_5[950];
    assign inter_6[951] = inter_5[951];
    assign inter_6[952] = inter_5[952];
    assign inter_6[953] = inter_5[953];
    assign inter_6[954] = inter_5[954];
    assign inter_6[955] = inter_5[955];
    assign inter_6[956] = inter_5[956];
    assign inter_6[957] = inter_5[957];
    assign inter_6[958] = inter_5[958];
    assign inter_6[959] = inter_5[959];
    assign inter_6[960] = inter_5[960]^inter_5[992];
    assign inter_6[961] = inter_5[961]^inter_5[993];
    assign inter_6[962] = inter_5[962]^inter_5[994];
    assign inter_6[963] = inter_5[963]^inter_5[995];
    assign inter_6[964] = inter_5[964]^inter_5[996];
    assign inter_6[965] = inter_5[965]^inter_5[997];
    assign inter_6[966] = inter_5[966]^inter_5[998];
    assign inter_6[967] = inter_5[967]^inter_5[999];
    assign inter_6[968] = inter_5[968]^inter_5[1000];
    assign inter_6[969] = inter_5[969]^inter_5[1001];
    assign inter_6[970] = inter_5[970]^inter_5[1002];
    assign inter_6[971] = inter_5[971]^inter_5[1003];
    assign inter_6[972] = inter_5[972]^inter_5[1004];
    assign inter_6[973] = inter_5[973]^inter_5[1005];
    assign inter_6[974] = inter_5[974]^inter_5[1006];
    assign inter_6[975] = inter_5[975]^inter_5[1007];
    assign inter_6[976] = inter_5[976]^inter_5[1008];
    assign inter_6[977] = inter_5[977]^inter_5[1009];
    assign inter_6[978] = inter_5[978]^inter_5[1010];
    assign inter_6[979] = inter_5[979]^inter_5[1011];
    assign inter_6[980] = inter_5[980]^inter_5[1012];
    assign inter_6[981] = inter_5[981]^inter_5[1013];
    assign inter_6[982] = inter_5[982]^inter_5[1014];
    assign inter_6[983] = inter_5[983]^inter_5[1015];
    assign inter_6[984] = inter_5[984]^inter_5[1016];
    assign inter_6[985] = inter_5[985]^inter_5[1017];
    assign inter_6[986] = inter_5[986]^inter_5[1018];
    assign inter_6[987] = inter_5[987]^inter_5[1019];
    assign inter_6[988] = inter_5[988]^inter_5[1020];
    assign inter_6[989] = inter_5[989]^inter_5[1021];
    assign inter_6[990] = inter_5[990]^inter_5[1022];
    assign inter_6[991] = inter_5[991]^inter_5[1023];
    assign inter_6[992] = inter_5[992];
    assign inter_6[993] = inter_5[993];
    assign inter_6[994] = inter_5[994];
    assign inter_6[995] = inter_5[995];
    assign inter_6[996] = inter_5[996];
    assign inter_6[997] = inter_5[997];
    assign inter_6[998] = inter_5[998];
    assign inter_6[999] = inter_5[999];
    assign inter_6[1000] = inter_5[1000];
    assign inter_6[1001] = inter_5[1001];
    assign inter_6[1002] = inter_5[1002];
    assign inter_6[1003] = inter_5[1003];
    assign inter_6[1004] = inter_5[1004];
    assign inter_6[1005] = inter_5[1005];
    assign inter_6[1006] = inter_5[1006];
    assign inter_6[1007] = inter_5[1007];
    assign inter_6[1008] = inter_5[1008];
    assign inter_6[1009] = inter_5[1009];
    assign inter_6[1010] = inter_5[1010];
    assign inter_6[1011] = inter_5[1011];
    assign inter_6[1012] = inter_5[1012];
    assign inter_6[1013] = inter_5[1013];
    assign inter_6[1014] = inter_5[1014];
    assign inter_6[1015] = inter_5[1015];
    assign inter_6[1016] = inter_5[1016];
    assign inter_6[1017] = inter_5[1017];
    assign inter_6[1018] = inter_5[1018];
    assign inter_6[1019] = inter_5[1019];
    assign inter_6[1020] = inter_5[1020];
    assign inter_6[1021] = inter_5[1021];
    assign inter_6[1022] = inter_5[1022];
    assign inter_6[1023] = inter_5[1023];
    /***************************/
    assign inter_7[0] = inter_6[0]^inter_6[64];
    assign inter_7[1] = inter_6[1]^inter_6[65];
    assign inter_7[2] = inter_6[2]^inter_6[66];
    assign inter_7[3] = inter_6[3]^inter_6[67];
    assign inter_7[4] = inter_6[4]^inter_6[68];
    assign inter_7[5] = inter_6[5]^inter_6[69];
    assign inter_7[6] = inter_6[6]^inter_6[70];
    assign inter_7[7] = inter_6[7]^inter_6[71];
    assign inter_7[8] = inter_6[8]^inter_6[72];
    assign inter_7[9] = inter_6[9]^inter_6[73];
    assign inter_7[10] = inter_6[10]^inter_6[74];
    assign inter_7[11] = inter_6[11]^inter_6[75];
    assign inter_7[12] = inter_6[12]^inter_6[76];
    assign inter_7[13] = inter_6[13]^inter_6[77];
    assign inter_7[14] = inter_6[14]^inter_6[78];
    assign inter_7[15] = inter_6[15]^inter_6[79];
    assign inter_7[16] = inter_6[16]^inter_6[80];
    assign inter_7[17] = inter_6[17]^inter_6[81];
    assign inter_7[18] = inter_6[18]^inter_6[82];
    assign inter_7[19] = inter_6[19]^inter_6[83];
    assign inter_7[20] = inter_6[20]^inter_6[84];
    assign inter_7[21] = inter_6[21]^inter_6[85];
    assign inter_7[22] = inter_6[22]^inter_6[86];
    assign inter_7[23] = inter_6[23]^inter_6[87];
    assign inter_7[24] = inter_6[24]^inter_6[88];
    assign inter_7[25] = inter_6[25]^inter_6[89];
    assign inter_7[26] = inter_6[26]^inter_6[90];
    assign inter_7[27] = inter_6[27]^inter_6[91];
    assign inter_7[28] = inter_6[28]^inter_6[92];
    assign inter_7[29] = inter_6[29]^inter_6[93];
    assign inter_7[30] = inter_6[30]^inter_6[94];
    assign inter_7[31] = inter_6[31]^inter_6[95];
    assign inter_7[32] = inter_6[32]^inter_6[96];
    assign inter_7[33] = inter_6[33]^inter_6[97];
    assign inter_7[34] = inter_6[34]^inter_6[98];
    assign inter_7[35] = inter_6[35]^inter_6[99];
    assign inter_7[36] = inter_6[36]^inter_6[100];
    assign inter_7[37] = inter_6[37]^inter_6[101];
    assign inter_7[38] = inter_6[38]^inter_6[102];
    assign inter_7[39] = inter_6[39]^inter_6[103];
    assign inter_7[40] = inter_6[40]^inter_6[104];
    assign inter_7[41] = inter_6[41]^inter_6[105];
    assign inter_7[42] = inter_6[42]^inter_6[106];
    assign inter_7[43] = inter_6[43]^inter_6[107];
    assign inter_7[44] = inter_6[44]^inter_6[108];
    assign inter_7[45] = inter_6[45]^inter_6[109];
    assign inter_7[46] = inter_6[46]^inter_6[110];
    assign inter_7[47] = inter_6[47]^inter_6[111];
    assign inter_7[48] = inter_6[48]^inter_6[112];
    assign inter_7[49] = inter_6[49]^inter_6[113];
    assign inter_7[50] = inter_6[50]^inter_6[114];
    assign inter_7[51] = inter_6[51]^inter_6[115];
    assign inter_7[52] = inter_6[52]^inter_6[116];
    assign inter_7[53] = inter_6[53]^inter_6[117];
    assign inter_7[54] = inter_6[54]^inter_6[118];
    assign inter_7[55] = inter_6[55]^inter_6[119];
    assign inter_7[56] = inter_6[56]^inter_6[120];
    assign inter_7[57] = inter_6[57]^inter_6[121];
    assign inter_7[58] = inter_6[58]^inter_6[122];
    assign inter_7[59] = inter_6[59]^inter_6[123];
    assign inter_7[60] = inter_6[60]^inter_6[124];
    assign inter_7[61] = inter_6[61]^inter_6[125];
    assign inter_7[62] = inter_6[62]^inter_6[126];
    assign inter_7[63] = inter_6[63]^inter_6[127];
    assign inter_7[64] = inter_6[64];
    assign inter_7[65] = inter_6[65];
    assign inter_7[66] = inter_6[66];
    assign inter_7[67] = inter_6[67];
    assign inter_7[68] = inter_6[68];
    assign inter_7[69] = inter_6[69];
    assign inter_7[70] = inter_6[70];
    assign inter_7[71] = inter_6[71];
    assign inter_7[72] = inter_6[72];
    assign inter_7[73] = inter_6[73];
    assign inter_7[74] = inter_6[74];
    assign inter_7[75] = inter_6[75];
    assign inter_7[76] = inter_6[76];
    assign inter_7[77] = inter_6[77];
    assign inter_7[78] = inter_6[78];
    assign inter_7[79] = inter_6[79];
    assign inter_7[80] = inter_6[80];
    assign inter_7[81] = inter_6[81];
    assign inter_7[82] = inter_6[82];
    assign inter_7[83] = inter_6[83];
    assign inter_7[84] = inter_6[84];
    assign inter_7[85] = inter_6[85];
    assign inter_7[86] = inter_6[86];
    assign inter_7[87] = inter_6[87];
    assign inter_7[88] = inter_6[88];
    assign inter_7[89] = inter_6[89];
    assign inter_7[90] = inter_6[90];
    assign inter_7[91] = inter_6[91];
    assign inter_7[92] = inter_6[92];
    assign inter_7[93] = inter_6[93];
    assign inter_7[94] = inter_6[94];
    assign inter_7[95] = inter_6[95];
    assign inter_7[96] = inter_6[96];
    assign inter_7[97] = inter_6[97];
    assign inter_7[98] = inter_6[98];
    assign inter_7[99] = inter_6[99];
    assign inter_7[100] = inter_6[100];
    assign inter_7[101] = inter_6[101];
    assign inter_7[102] = inter_6[102];
    assign inter_7[103] = inter_6[103];
    assign inter_7[104] = inter_6[104];
    assign inter_7[105] = inter_6[105];
    assign inter_7[106] = inter_6[106];
    assign inter_7[107] = inter_6[107];
    assign inter_7[108] = inter_6[108];
    assign inter_7[109] = inter_6[109];
    assign inter_7[110] = inter_6[110];
    assign inter_7[111] = inter_6[111];
    assign inter_7[112] = inter_6[112];
    assign inter_7[113] = inter_6[113];
    assign inter_7[114] = inter_6[114];
    assign inter_7[115] = inter_6[115];
    assign inter_7[116] = inter_6[116];
    assign inter_7[117] = inter_6[117];
    assign inter_7[118] = inter_6[118];
    assign inter_7[119] = inter_6[119];
    assign inter_7[120] = inter_6[120];
    assign inter_7[121] = inter_6[121];
    assign inter_7[122] = inter_6[122];
    assign inter_7[123] = inter_6[123];
    assign inter_7[124] = inter_6[124];
    assign inter_7[125] = inter_6[125];
    assign inter_7[126] = inter_6[126];
    assign inter_7[127] = inter_6[127];
    assign inter_7[128] = inter_6[128]^inter_6[192];
    assign inter_7[129] = inter_6[129]^inter_6[193];
    assign inter_7[130] = inter_6[130]^inter_6[194];
    assign inter_7[131] = inter_6[131]^inter_6[195];
    assign inter_7[132] = inter_6[132]^inter_6[196];
    assign inter_7[133] = inter_6[133]^inter_6[197];
    assign inter_7[134] = inter_6[134]^inter_6[198];
    assign inter_7[135] = inter_6[135]^inter_6[199];
    assign inter_7[136] = inter_6[136]^inter_6[200];
    assign inter_7[137] = inter_6[137]^inter_6[201];
    assign inter_7[138] = inter_6[138]^inter_6[202];
    assign inter_7[139] = inter_6[139]^inter_6[203];
    assign inter_7[140] = inter_6[140]^inter_6[204];
    assign inter_7[141] = inter_6[141]^inter_6[205];
    assign inter_7[142] = inter_6[142]^inter_6[206];
    assign inter_7[143] = inter_6[143]^inter_6[207];
    assign inter_7[144] = inter_6[144]^inter_6[208];
    assign inter_7[145] = inter_6[145]^inter_6[209];
    assign inter_7[146] = inter_6[146]^inter_6[210];
    assign inter_7[147] = inter_6[147]^inter_6[211];
    assign inter_7[148] = inter_6[148]^inter_6[212];
    assign inter_7[149] = inter_6[149]^inter_6[213];
    assign inter_7[150] = inter_6[150]^inter_6[214];
    assign inter_7[151] = inter_6[151]^inter_6[215];
    assign inter_7[152] = inter_6[152]^inter_6[216];
    assign inter_7[153] = inter_6[153]^inter_6[217];
    assign inter_7[154] = inter_6[154]^inter_6[218];
    assign inter_7[155] = inter_6[155]^inter_6[219];
    assign inter_7[156] = inter_6[156]^inter_6[220];
    assign inter_7[157] = inter_6[157]^inter_6[221];
    assign inter_7[158] = inter_6[158]^inter_6[222];
    assign inter_7[159] = inter_6[159]^inter_6[223];
    assign inter_7[160] = inter_6[160]^inter_6[224];
    assign inter_7[161] = inter_6[161]^inter_6[225];
    assign inter_7[162] = inter_6[162]^inter_6[226];
    assign inter_7[163] = inter_6[163]^inter_6[227];
    assign inter_7[164] = inter_6[164]^inter_6[228];
    assign inter_7[165] = inter_6[165]^inter_6[229];
    assign inter_7[166] = inter_6[166]^inter_6[230];
    assign inter_7[167] = inter_6[167]^inter_6[231];
    assign inter_7[168] = inter_6[168]^inter_6[232];
    assign inter_7[169] = inter_6[169]^inter_6[233];
    assign inter_7[170] = inter_6[170]^inter_6[234];
    assign inter_7[171] = inter_6[171]^inter_6[235];
    assign inter_7[172] = inter_6[172]^inter_6[236];
    assign inter_7[173] = inter_6[173]^inter_6[237];
    assign inter_7[174] = inter_6[174]^inter_6[238];
    assign inter_7[175] = inter_6[175]^inter_6[239];
    assign inter_7[176] = inter_6[176]^inter_6[240];
    assign inter_7[177] = inter_6[177]^inter_6[241];
    assign inter_7[178] = inter_6[178]^inter_6[242];
    assign inter_7[179] = inter_6[179]^inter_6[243];
    assign inter_7[180] = inter_6[180]^inter_6[244];
    assign inter_7[181] = inter_6[181]^inter_6[245];
    assign inter_7[182] = inter_6[182]^inter_6[246];
    assign inter_7[183] = inter_6[183]^inter_6[247];
    assign inter_7[184] = inter_6[184]^inter_6[248];
    assign inter_7[185] = inter_6[185]^inter_6[249];
    assign inter_7[186] = inter_6[186]^inter_6[250];
    assign inter_7[187] = inter_6[187]^inter_6[251];
    assign inter_7[188] = inter_6[188]^inter_6[252];
    assign inter_7[189] = inter_6[189]^inter_6[253];
    assign inter_7[190] = inter_6[190]^inter_6[254];
    assign inter_7[191] = inter_6[191]^inter_6[255];
    assign inter_7[192] = inter_6[192];
    assign inter_7[193] = inter_6[193];
    assign inter_7[194] = inter_6[194];
    assign inter_7[195] = inter_6[195];
    assign inter_7[196] = inter_6[196];
    assign inter_7[197] = inter_6[197];
    assign inter_7[198] = inter_6[198];
    assign inter_7[199] = inter_6[199];
    assign inter_7[200] = inter_6[200];
    assign inter_7[201] = inter_6[201];
    assign inter_7[202] = inter_6[202];
    assign inter_7[203] = inter_6[203];
    assign inter_7[204] = inter_6[204];
    assign inter_7[205] = inter_6[205];
    assign inter_7[206] = inter_6[206];
    assign inter_7[207] = inter_6[207];
    assign inter_7[208] = inter_6[208];
    assign inter_7[209] = inter_6[209];
    assign inter_7[210] = inter_6[210];
    assign inter_7[211] = inter_6[211];
    assign inter_7[212] = inter_6[212];
    assign inter_7[213] = inter_6[213];
    assign inter_7[214] = inter_6[214];
    assign inter_7[215] = inter_6[215];
    assign inter_7[216] = inter_6[216];
    assign inter_7[217] = inter_6[217];
    assign inter_7[218] = inter_6[218];
    assign inter_7[219] = inter_6[219];
    assign inter_7[220] = inter_6[220];
    assign inter_7[221] = inter_6[221];
    assign inter_7[222] = inter_6[222];
    assign inter_7[223] = inter_6[223];
    assign inter_7[224] = inter_6[224];
    assign inter_7[225] = inter_6[225];
    assign inter_7[226] = inter_6[226];
    assign inter_7[227] = inter_6[227];
    assign inter_7[228] = inter_6[228];
    assign inter_7[229] = inter_6[229];
    assign inter_7[230] = inter_6[230];
    assign inter_7[231] = inter_6[231];
    assign inter_7[232] = inter_6[232];
    assign inter_7[233] = inter_6[233];
    assign inter_7[234] = inter_6[234];
    assign inter_7[235] = inter_6[235];
    assign inter_7[236] = inter_6[236];
    assign inter_7[237] = inter_6[237];
    assign inter_7[238] = inter_6[238];
    assign inter_7[239] = inter_6[239];
    assign inter_7[240] = inter_6[240];
    assign inter_7[241] = inter_6[241];
    assign inter_7[242] = inter_6[242];
    assign inter_7[243] = inter_6[243];
    assign inter_7[244] = inter_6[244];
    assign inter_7[245] = inter_6[245];
    assign inter_7[246] = inter_6[246];
    assign inter_7[247] = inter_6[247];
    assign inter_7[248] = inter_6[248];
    assign inter_7[249] = inter_6[249];
    assign inter_7[250] = inter_6[250];
    assign inter_7[251] = inter_6[251];
    assign inter_7[252] = inter_6[252];
    assign inter_7[253] = inter_6[253];
    assign inter_7[254] = inter_6[254];
    assign inter_7[255] = inter_6[255];
    assign inter_7[256] = inter_6[256]^inter_6[320];
    assign inter_7[257] = inter_6[257]^inter_6[321];
    assign inter_7[258] = inter_6[258]^inter_6[322];
    assign inter_7[259] = inter_6[259]^inter_6[323];
    assign inter_7[260] = inter_6[260]^inter_6[324];
    assign inter_7[261] = inter_6[261]^inter_6[325];
    assign inter_7[262] = inter_6[262]^inter_6[326];
    assign inter_7[263] = inter_6[263]^inter_6[327];
    assign inter_7[264] = inter_6[264]^inter_6[328];
    assign inter_7[265] = inter_6[265]^inter_6[329];
    assign inter_7[266] = inter_6[266]^inter_6[330];
    assign inter_7[267] = inter_6[267]^inter_6[331];
    assign inter_7[268] = inter_6[268]^inter_6[332];
    assign inter_7[269] = inter_6[269]^inter_6[333];
    assign inter_7[270] = inter_6[270]^inter_6[334];
    assign inter_7[271] = inter_6[271]^inter_6[335];
    assign inter_7[272] = inter_6[272]^inter_6[336];
    assign inter_7[273] = inter_6[273]^inter_6[337];
    assign inter_7[274] = inter_6[274]^inter_6[338];
    assign inter_7[275] = inter_6[275]^inter_6[339];
    assign inter_7[276] = inter_6[276]^inter_6[340];
    assign inter_7[277] = inter_6[277]^inter_6[341];
    assign inter_7[278] = inter_6[278]^inter_6[342];
    assign inter_7[279] = inter_6[279]^inter_6[343];
    assign inter_7[280] = inter_6[280]^inter_6[344];
    assign inter_7[281] = inter_6[281]^inter_6[345];
    assign inter_7[282] = inter_6[282]^inter_6[346];
    assign inter_7[283] = inter_6[283]^inter_6[347];
    assign inter_7[284] = inter_6[284]^inter_6[348];
    assign inter_7[285] = inter_6[285]^inter_6[349];
    assign inter_7[286] = inter_6[286]^inter_6[350];
    assign inter_7[287] = inter_6[287]^inter_6[351];
    assign inter_7[288] = inter_6[288]^inter_6[352];
    assign inter_7[289] = inter_6[289]^inter_6[353];
    assign inter_7[290] = inter_6[290]^inter_6[354];
    assign inter_7[291] = inter_6[291]^inter_6[355];
    assign inter_7[292] = inter_6[292]^inter_6[356];
    assign inter_7[293] = inter_6[293]^inter_6[357];
    assign inter_7[294] = inter_6[294]^inter_6[358];
    assign inter_7[295] = inter_6[295]^inter_6[359];
    assign inter_7[296] = inter_6[296]^inter_6[360];
    assign inter_7[297] = inter_6[297]^inter_6[361];
    assign inter_7[298] = inter_6[298]^inter_6[362];
    assign inter_7[299] = inter_6[299]^inter_6[363];
    assign inter_7[300] = inter_6[300]^inter_6[364];
    assign inter_7[301] = inter_6[301]^inter_6[365];
    assign inter_7[302] = inter_6[302]^inter_6[366];
    assign inter_7[303] = inter_6[303]^inter_6[367];
    assign inter_7[304] = inter_6[304]^inter_6[368];
    assign inter_7[305] = inter_6[305]^inter_6[369];
    assign inter_7[306] = inter_6[306]^inter_6[370];
    assign inter_7[307] = inter_6[307]^inter_6[371];
    assign inter_7[308] = inter_6[308]^inter_6[372];
    assign inter_7[309] = inter_6[309]^inter_6[373];
    assign inter_7[310] = inter_6[310]^inter_6[374];
    assign inter_7[311] = inter_6[311]^inter_6[375];
    assign inter_7[312] = inter_6[312]^inter_6[376];
    assign inter_7[313] = inter_6[313]^inter_6[377];
    assign inter_7[314] = inter_6[314]^inter_6[378];
    assign inter_7[315] = inter_6[315]^inter_6[379];
    assign inter_7[316] = inter_6[316]^inter_6[380];
    assign inter_7[317] = inter_6[317]^inter_6[381];
    assign inter_7[318] = inter_6[318]^inter_6[382];
    assign inter_7[319] = inter_6[319]^inter_6[383];
    assign inter_7[320] = inter_6[320];
    assign inter_7[321] = inter_6[321];
    assign inter_7[322] = inter_6[322];
    assign inter_7[323] = inter_6[323];
    assign inter_7[324] = inter_6[324];
    assign inter_7[325] = inter_6[325];
    assign inter_7[326] = inter_6[326];
    assign inter_7[327] = inter_6[327];
    assign inter_7[328] = inter_6[328];
    assign inter_7[329] = inter_6[329];
    assign inter_7[330] = inter_6[330];
    assign inter_7[331] = inter_6[331];
    assign inter_7[332] = inter_6[332];
    assign inter_7[333] = inter_6[333];
    assign inter_7[334] = inter_6[334];
    assign inter_7[335] = inter_6[335];
    assign inter_7[336] = inter_6[336];
    assign inter_7[337] = inter_6[337];
    assign inter_7[338] = inter_6[338];
    assign inter_7[339] = inter_6[339];
    assign inter_7[340] = inter_6[340];
    assign inter_7[341] = inter_6[341];
    assign inter_7[342] = inter_6[342];
    assign inter_7[343] = inter_6[343];
    assign inter_7[344] = inter_6[344];
    assign inter_7[345] = inter_6[345];
    assign inter_7[346] = inter_6[346];
    assign inter_7[347] = inter_6[347];
    assign inter_7[348] = inter_6[348];
    assign inter_7[349] = inter_6[349];
    assign inter_7[350] = inter_6[350];
    assign inter_7[351] = inter_6[351];
    assign inter_7[352] = inter_6[352];
    assign inter_7[353] = inter_6[353];
    assign inter_7[354] = inter_6[354];
    assign inter_7[355] = inter_6[355];
    assign inter_7[356] = inter_6[356];
    assign inter_7[357] = inter_6[357];
    assign inter_7[358] = inter_6[358];
    assign inter_7[359] = inter_6[359];
    assign inter_7[360] = inter_6[360];
    assign inter_7[361] = inter_6[361];
    assign inter_7[362] = inter_6[362];
    assign inter_7[363] = inter_6[363];
    assign inter_7[364] = inter_6[364];
    assign inter_7[365] = inter_6[365];
    assign inter_7[366] = inter_6[366];
    assign inter_7[367] = inter_6[367];
    assign inter_7[368] = inter_6[368];
    assign inter_7[369] = inter_6[369];
    assign inter_7[370] = inter_6[370];
    assign inter_7[371] = inter_6[371];
    assign inter_7[372] = inter_6[372];
    assign inter_7[373] = inter_6[373];
    assign inter_7[374] = inter_6[374];
    assign inter_7[375] = inter_6[375];
    assign inter_7[376] = inter_6[376];
    assign inter_7[377] = inter_6[377];
    assign inter_7[378] = inter_6[378];
    assign inter_7[379] = inter_6[379];
    assign inter_7[380] = inter_6[380];
    assign inter_7[381] = inter_6[381];
    assign inter_7[382] = inter_6[382];
    assign inter_7[383] = inter_6[383];
    assign inter_7[384] = inter_6[384]^inter_6[448];
    assign inter_7[385] = inter_6[385]^inter_6[449];
    assign inter_7[386] = inter_6[386]^inter_6[450];
    assign inter_7[387] = inter_6[387]^inter_6[451];
    assign inter_7[388] = inter_6[388]^inter_6[452];
    assign inter_7[389] = inter_6[389]^inter_6[453];
    assign inter_7[390] = inter_6[390]^inter_6[454];
    assign inter_7[391] = inter_6[391]^inter_6[455];
    assign inter_7[392] = inter_6[392]^inter_6[456];
    assign inter_7[393] = inter_6[393]^inter_6[457];
    assign inter_7[394] = inter_6[394]^inter_6[458];
    assign inter_7[395] = inter_6[395]^inter_6[459];
    assign inter_7[396] = inter_6[396]^inter_6[460];
    assign inter_7[397] = inter_6[397]^inter_6[461];
    assign inter_7[398] = inter_6[398]^inter_6[462];
    assign inter_7[399] = inter_6[399]^inter_6[463];
    assign inter_7[400] = inter_6[400]^inter_6[464];
    assign inter_7[401] = inter_6[401]^inter_6[465];
    assign inter_7[402] = inter_6[402]^inter_6[466];
    assign inter_7[403] = inter_6[403]^inter_6[467];
    assign inter_7[404] = inter_6[404]^inter_6[468];
    assign inter_7[405] = inter_6[405]^inter_6[469];
    assign inter_7[406] = inter_6[406]^inter_6[470];
    assign inter_7[407] = inter_6[407]^inter_6[471];
    assign inter_7[408] = inter_6[408]^inter_6[472];
    assign inter_7[409] = inter_6[409]^inter_6[473];
    assign inter_7[410] = inter_6[410]^inter_6[474];
    assign inter_7[411] = inter_6[411]^inter_6[475];
    assign inter_7[412] = inter_6[412]^inter_6[476];
    assign inter_7[413] = inter_6[413]^inter_6[477];
    assign inter_7[414] = inter_6[414]^inter_6[478];
    assign inter_7[415] = inter_6[415]^inter_6[479];
    assign inter_7[416] = inter_6[416]^inter_6[480];
    assign inter_7[417] = inter_6[417]^inter_6[481];
    assign inter_7[418] = inter_6[418]^inter_6[482];
    assign inter_7[419] = inter_6[419]^inter_6[483];
    assign inter_7[420] = inter_6[420]^inter_6[484];
    assign inter_7[421] = inter_6[421]^inter_6[485];
    assign inter_7[422] = inter_6[422]^inter_6[486];
    assign inter_7[423] = inter_6[423]^inter_6[487];
    assign inter_7[424] = inter_6[424]^inter_6[488];
    assign inter_7[425] = inter_6[425]^inter_6[489];
    assign inter_7[426] = inter_6[426]^inter_6[490];
    assign inter_7[427] = inter_6[427]^inter_6[491];
    assign inter_7[428] = inter_6[428]^inter_6[492];
    assign inter_7[429] = inter_6[429]^inter_6[493];
    assign inter_7[430] = inter_6[430]^inter_6[494];
    assign inter_7[431] = inter_6[431]^inter_6[495];
    assign inter_7[432] = inter_6[432]^inter_6[496];
    assign inter_7[433] = inter_6[433]^inter_6[497];
    assign inter_7[434] = inter_6[434]^inter_6[498];
    assign inter_7[435] = inter_6[435]^inter_6[499];
    assign inter_7[436] = inter_6[436]^inter_6[500];
    assign inter_7[437] = inter_6[437]^inter_6[501];
    assign inter_7[438] = inter_6[438]^inter_6[502];
    assign inter_7[439] = inter_6[439]^inter_6[503];
    assign inter_7[440] = inter_6[440]^inter_6[504];
    assign inter_7[441] = inter_6[441]^inter_6[505];
    assign inter_7[442] = inter_6[442]^inter_6[506];
    assign inter_7[443] = inter_6[443]^inter_6[507];
    assign inter_7[444] = inter_6[444]^inter_6[508];
    assign inter_7[445] = inter_6[445]^inter_6[509];
    assign inter_7[446] = inter_6[446]^inter_6[510];
    assign inter_7[447] = inter_6[447]^inter_6[511];
    assign inter_7[448] = inter_6[448];
    assign inter_7[449] = inter_6[449];
    assign inter_7[450] = inter_6[450];
    assign inter_7[451] = inter_6[451];
    assign inter_7[452] = inter_6[452];
    assign inter_7[453] = inter_6[453];
    assign inter_7[454] = inter_6[454];
    assign inter_7[455] = inter_6[455];
    assign inter_7[456] = inter_6[456];
    assign inter_7[457] = inter_6[457];
    assign inter_7[458] = inter_6[458];
    assign inter_7[459] = inter_6[459];
    assign inter_7[460] = inter_6[460];
    assign inter_7[461] = inter_6[461];
    assign inter_7[462] = inter_6[462];
    assign inter_7[463] = inter_6[463];
    assign inter_7[464] = inter_6[464];
    assign inter_7[465] = inter_6[465];
    assign inter_7[466] = inter_6[466];
    assign inter_7[467] = inter_6[467];
    assign inter_7[468] = inter_6[468];
    assign inter_7[469] = inter_6[469];
    assign inter_7[470] = inter_6[470];
    assign inter_7[471] = inter_6[471];
    assign inter_7[472] = inter_6[472];
    assign inter_7[473] = inter_6[473];
    assign inter_7[474] = inter_6[474];
    assign inter_7[475] = inter_6[475];
    assign inter_7[476] = inter_6[476];
    assign inter_7[477] = inter_6[477];
    assign inter_7[478] = inter_6[478];
    assign inter_7[479] = inter_6[479];
    assign inter_7[480] = inter_6[480];
    assign inter_7[481] = inter_6[481];
    assign inter_7[482] = inter_6[482];
    assign inter_7[483] = inter_6[483];
    assign inter_7[484] = inter_6[484];
    assign inter_7[485] = inter_6[485];
    assign inter_7[486] = inter_6[486];
    assign inter_7[487] = inter_6[487];
    assign inter_7[488] = inter_6[488];
    assign inter_7[489] = inter_6[489];
    assign inter_7[490] = inter_6[490];
    assign inter_7[491] = inter_6[491];
    assign inter_7[492] = inter_6[492];
    assign inter_7[493] = inter_6[493];
    assign inter_7[494] = inter_6[494];
    assign inter_7[495] = inter_6[495];
    assign inter_7[496] = inter_6[496];
    assign inter_7[497] = inter_6[497];
    assign inter_7[498] = inter_6[498];
    assign inter_7[499] = inter_6[499];
    assign inter_7[500] = inter_6[500];
    assign inter_7[501] = inter_6[501];
    assign inter_7[502] = inter_6[502];
    assign inter_7[503] = inter_6[503];
    assign inter_7[504] = inter_6[504];
    assign inter_7[505] = inter_6[505];
    assign inter_7[506] = inter_6[506];
    assign inter_7[507] = inter_6[507];
    assign inter_7[508] = inter_6[508];
    assign inter_7[509] = inter_6[509];
    assign inter_7[510] = inter_6[510];
    assign inter_7[511] = inter_6[511];
    assign inter_7[512] = inter_6[512]^inter_6[576];
    assign inter_7[513] = inter_6[513]^inter_6[577];
    assign inter_7[514] = inter_6[514]^inter_6[578];
    assign inter_7[515] = inter_6[515]^inter_6[579];
    assign inter_7[516] = inter_6[516]^inter_6[580];
    assign inter_7[517] = inter_6[517]^inter_6[581];
    assign inter_7[518] = inter_6[518]^inter_6[582];
    assign inter_7[519] = inter_6[519]^inter_6[583];
    assign inter_7[520] = inter_6[520]^inter_6[584];
    assign inter_7[521] = inter_6[521]^inter_6[585];
    assign inter_7[522] = inter_6[522]^inter_6[586];
    assign inter_7[523] = inter_6[523]^inter_6[587];
    assign inter_7[524] = inter_6[524]^inter_6[588];
    assign inter_7[525] = inter_6[525]^inter_6[589];
    assign inter_7[526] = inter_6[526]^inter_6[590];
    assign inter_7[527] = inter_6[527]^inter_6[591];
    assign inter_7[528] = inter_6[528]^inter_6[592];
    assign inter_7[529] = inter_6[529]^inter_6[593];
    assign inter_7[530] = inter_6[530]^inter_6[594];
    assign inter_7[531] = inter_6[531]^inter_6[595];
    assign inter_7[532] = inter_6[532]^inter_6[596];
    assign inter_7[533] = inter_6[533]^inter_6[597];
    assign inter_7[534] = inter_6[534]^inter_6[598];
    assign inter_7[535] = inter_6[535]^inter_6[599];
    assign inter_7[536] = inter_6[536]^inter_6[600];
    assign inter_7[537] = inter_6[537]^inter_6[601];
    assign inter_7[538] = inter_6[538]^inter_6[602];
    assign inter_7[539] = inter_6[539]^inter_6[603];
    assign inter_7[540] = inter_6[540]^inter_6[604];
    assign inter_7[541] = inter_6[541]^inter_6[605];
    assign inter_7[542] = inter_6[542]^inter_6[606];
    assign inter_7[543] = inter_6[543]^inter_6[607];
    assign inter_7[544] = inter_6[544]^inter_6[608];
    assign inter_7[545] = inter_6[545]^inter_6[609];
    assign inter_7[546] = inter_6[546]^inter_6[610];
    assign inter_7[547] = inter_6[547]^inter_6[611];
    assign inter_7[548] = inter_6[548]^inter_6[612];
    assign inter_7[549] = inter_6[549]^inter_6[613];
    assign inter_7[550] = inter_6[550]^inter_6[614];
    assign inter_7[551] = inter_6[551]^inter_6[615];
    assign inter_7[552] = inter_6[552]^inter_6[616];
    assign inter_7[553] = inter_6[553]^inter_6[617];
    assign inter_7[554] = inter_6[554]^inter_6[618];
    assign inter_7[555] = inter_6[555]^inter_6[619];
    assign inter_7[556] = inter_6[556]^inter_6[620];
    assign inter_7[557] = inter_6[557]^inter_6[621];
    assign inter_7[558] = inter_6[558]^inter_6[622];
    assign inter_7[559] = inter_6[559]^inter_6[623];
    assign inter_7[560] = inter_6[560]^inter_6[624];
    assign inter_7[561] = inter_6[561]^inter_6[625];
    assign inter_7[562] = inter_6[562]^inter_6[626];
    assign inter_7[563] = inter_6[563]^inter_6[627];
    assign inter_7[564] = inter_6[564]^inter_6[628];
    assign inter_7[565] = inter_6[565]^inter_6[629];
    assign inter_7[566] = inter_6[566]^inter_6[630];
    assign inter_7[567] = inter_6[567]^inter_6[631];
    assign inter_7[568] = inter_6[568]^inter_6[632];
    assign inter_7[569] = inter_6[569]^inter_6[633];
    assign inter_7[570] = inter_6[570]^inter_6[634];
    assign inter_7[571] = inter_6[571]^inter_6[635];
    assign inter_7[572] = inter_6[572]^inter_6[636];
    assign inter_7[573] = inter_6[573]^inter_6[637];
    assign inter_7[574] = inter_6[574]^inter_6[638];
    assign inter_7[575] = inter_6[575]^inter_6[639];
    assign inter_7[576] = inter_6[576];
    assign inter_7[577] = inter_6[577];
    assign inter_7[578] = inter_6[578];
    assign inter_7[579] = inter_6[579];
    assign inter_7[580] = inter_6[580];
    assign inter_7[581] = inter_6[581];
    assign inter_7[582] = inter_6[582];
    assign inter_7[583] = inter_6[583];
    assign inter_7[584] = inter_6[584];
    assign inter_7[585] = inter_6[585];
    assign inter_7[586] = inter_6[586];
    assign inter_7[587] = inter_6[587];
    assign inter_7[588] = inter_6[588];
    assign inter_7[589] = inter_6[589];
    assign inter_7[590] = inter_6[590];
    assign inter_7[591] = inter_6[591];
    assign inter_7[592] = inter_6[592];
    assign inter_7[593] = inter_6[593];
    assign inter_7[594] = inter_6[594];
    assign inter_7[595] = inter_6[595];
    assign inter_7[596] = inter_6[596];
    assign inter_7[597] = inter_6[597];
    assign inter_7[598] = inter_6[598];
    assign inter_7[599] = inter_6[599];
    assign inter_7[600] = inter_6[600];
    assign inter_7[601] = inter_6[601];
    assign inter_7[602] = inter_6[602];
    assign inter_7[603] = inter_6[603];
    assign inter_7[604] = inter_6[604];
    assign inter_7[605] = inter_6[605];
    assign inter_7[606] = inter_6[606];
    assign inter_7[607] = inter_6[607];
    assign inter_7[608] = inter_6[608];
    assign inter_7[609] = inter_6[609];
    assign inter_7[610] = inter_6[610];
    assign inter_7[611] = inter_6[611];
    assign inter_7[612] = inter_6[612];
    assign inter_7[613] = inter_6[613];
    assign inter_7[614] = inter_6[614];
    assign inter_7[615] = inter_6[615];
    assign inter_7[616] = inter_6[616];
    assign inter_7[617] = inter_6[617];
    assign inter_7[618] = inter_6[618];
    assign inter_7[619] = inter_6[619];
    assign inter_7[620] = inter_6[620];
    assign inter_7[621] = inter_6[621];
    assign inter_7[622] = inter_6[622];
    assign inter_7[623] = inter_6[623];
    assign inter_7[624] = inter_6[624];
    assign inter_7[625] = inter_6[625];
    assign inter_7[626] = inter_6[626];
    assign inter_7[627] = inter_6[627];
    assign inter_7[628] = inter_6[628];
    assign inter_7[629] = inter_6[629];
    assign inter_7[630] = inter_6[630];
    assign inter_7[631] = inter_6[631];
    assign inter_7[632] = inter_6[632];
    assign inter_7[633] = inter_6[633];
    assign inter_7[634] = inter_6[634];
    assign inter_7[635] = inter_6[635];
    assign inter_7[636] = inter_6[636];
    assign inter_7[637] = inter_6[637];
    assign inter_7[638] = inter_6[638];
    assign inter_7[639] = inter_6[639];
    assign inter_7[640] = inter_6[640]^inter_6[704];
    assign inter_7[641] = inter_6[641]^inter_6[705];
    assign inter_7[642] = inter_6[642]^inter_6[706];
    assign inter_7[643] = inter_6[643]^inter_6[707];
    assign inter_7[644] = inter_6[644]^inter_6[708];
    assign inter_7[645] = inter_6[645]^inter_6[709];
    assign inter_7[646] = inter_6[646]^inter_6[710];
    assign inter_7[647] = inter_6[647]^inter_6[711];
    assign inter_7[648] = inter_6[648]^inter_6[712];
    assign inter_7[649] = inter_6[649]^inter_6[713];
    assign inter_7[650] = inter_6[650]^inter_6[714];
    assign inter_7[651] = inter_6[651]^inter_6[715];
    assign inter_7[652] = inter_6[652]^inter_6[716];
    assign inter_7[653] = inter_6[653]^inter_6[717];
    assign inter_7[654] = inter_6[654]^inter_6[718];
    assign inter_7[655] = inter_6[655]^inter_6[719];
    assign inter_7[656] = inter_6[656]^inter_6[720];
    assign inter_7[657] = inter_6[657]^inter_6[721];
    assign inter_7[658] = inter_6[658]^inter_6[722];
    assign inter_7[659] = inter_6[659]^inter_6[723];
    assign inter_7[660] = inter_6[660]^inter_6[724];
    assign inter_7[661] = inter_6[661]^inter_6[725];
    assign inter_7[662] = inter_6[662]^inter_6[726];
    assign inter_7[663] = inter_6[663]^inter_6[727];
    assign inter_7[664] = inter_6[664]^inter_6[728];
    assign inter_7[665] = inter_6[665]^inter_6[729];
    assign inter_7[666] = inter_6[666]^inter_6[730];
    assign inter_7[667] = inter_6[667]^inter_6[731];
    assign inter_7[668] = inter_6[668]^inter_6[732];
    assign inter_7[669] = inter_6[669]^inter_6[733];
    assign inter_7[670] = inter_6[670]^inter_6[734];
    assign inter_7[671] = inter_6[671]^inter_6[735];
    assign inter_7[672] = inter_6[672]^inter_6[736];
    assign inter_7[673] = inter_6[673]^inter_6[737];
    assign inter_7[674] = inter_6[674]^inter_6[738];
    assign inter_7[675] = inter_6[675]^inter_6[739];
    assign inter_7[676] = inter_6[676]^inter_6[740];
    assign inter_7[677] = inter_6[677]^inter_6[741];
    assign inter_7[678] = inter_6[678]^inter_6[742];
    assign inter_7[679] = inter_6[679]^inter_6[743];
    assign inter_7[680] = inter_6[680]^inter_6[744];
    assign inter_7[681] = inter_6[681]^inter_6[745];
    assign inter_7[682] = inter_6[682]^inter_6[746];
    assign inter_7[683] = inter_6[683]^inter_6[747];
    assign inter_7[684] = inter_6[684]^inter_6[748];
    assign inter_7[685] = inter_6[685]^inter_6[749];
    assign inter_7[686] = inter_6[686]^inter_6[750];
    assign inter_7[687] = inter_6[687]^inter_6[751];
    assign inter_7[688] = inter_6[688]^inter_6[752];
    assign inter_7[689] = inter_6[689]^inter_6[753];
    assign inter_7[690] = inter_6[690]^inter_6[754];
    assign inter_7[691] = inter_6[691]^inter_6[755];
    assign inter_7[692] = inter_6[692]^inter_6[756];
    assign inter_7[693] = inter_6[693]^inter_6[757];
    assign inter_7[694] = inter_6[694]^inter_6[758];
    assign inter_7[695] = inter_6[695]^inter_6[759];
    assign inter_7[696] = inter_6[696]^inter_6[760];
    assign inter_7[697] = inter_6[697]^inter_6[761];
    assign inter_7[698] = inter_6[698]^inter_6[762];
    assign inter_7[699] = inter_6[699]^inter_6[763];
    assign inter_7[700] = inter_6[700]^inter_6[764];
    assign inter_7[701] = inter_6[701]^inter_6[765];
    assign inter_7[702] = inter_6[702]^inter_6[766];
    assign inter_7[703] = inter_6[703]^inter_6[767];
    assign inter_7[704] = inter_6[704];
    assign inter_7[705] = inter_6[705];
    assign inter_7[706] = inter_6[706];
    assign inter_7[707] = inter_6[707];
    assign inter_7[708] = inter_6[708];
    assign inter_7[709] = inter_6[709];
    assign inter_7[710] = inter_6[710];
    assign inter_7[711] = inter_6[711];
    assign inter_7[712] = inter_6[712];
    assign inter_7[713] = inter_6[713];
    assign inter_7[714] = inter_6[714];
    assign inter_7[715] = inter_6[715];
    assign inter_7[716] = inter_6[716];
    assign inter_7[717] = inter_6[717];
    assign inter_7[718] = inter_6[718];
    assign inter_7[719] = inter_6[719];
    assign inter_7[720] = inter_6[720];
    assign inter_7[721] = inter_6[721];
    assign inter_7[722] = inter_6[722];
    assign inter_7[723] = inter_6[723];
    assign inter_7[724] = inter_6[724];
    assign inter_7[725] = inter_6[725];
    assign inter_7[726] = inter_6[726];
    assign inter_7[727] = inter_6[727];
    assign inter_7[728] = inter_6[728];
    assign inter_7[729] = inter_6[729];
    assign inter_7[730] = inter_6[730];
    assign inter_7[731] = inter_6[731];
    assign inter_7[732] = inter_6[732];
    assign inter_7[733] = inter_6[733];
    assign inter_7[734] = inter_6[734];
    assign inter_7[735] = inter_6[735];
    assign inter_7[736] = inter_6[736];
    assign inter_7[737] = inter_6[737];
    assign inter_7[738] = inter_6[738];
    assign inter_7[739] = inter_6[739];
    assign inter_7[740] = inter_6[740];
    assign inter_7[741] = inter_6[741];
    assign inter_7[742] = inter_6[742];
    assign inter_7[743] = inter_6[743];
    assign inter_7[744] = inter_6[744];
    assign inter_7[745] = inter_6[745];
    assign inter_7[746] = inter_6[746];
    assign inter_7[747] = inter_6[747];
    assign inter_7[748] = inter_6[748];
    assign inter_7[749] = inter_6[749];
    assign inter_7[750] = inter_6[750];
    assign inter_7[751] = inter_6[751];
    assign inter_7[752] = inter_6[752];
    assign inter_7[753] = inter_6[753];
    assign inter_7[754] = inter_6[754];
    assign inter_7[755] = inter_6[755];
    assign inter_7[756] = inter_6[756];
    assign inter_7[757] = inter_6[757];
    assign inter_7[758] = inter_6[758];
    assign inter_7[759] = inter_6[759];
    assign inter_7[760] = inter_6[760];
    assign inter_7[761] = inter_6[761];
    assign inter_7[762] = inter_6[762];
    assign inter_7[763] = inter_6[763];
    assign inter_7[764] = inter_6[764];
    assign inter_7[765] = inter_6[765];
    assign inter_7[766] = inter_6[766];
    assign inter_7[767] = inter_6[767];
    assign inter_7[768] = inter_6[768]^inter_6[832];
    assign inter_7[769] = inter_6[769]^inter_6[833];
    assign inter_7[770] = inter_6[770]^inter_6[834];
    assign inter_7[771] = inter_6[771]^inter_6[835];
    assign inter_7[772] = inter_6[772]^inter_6[836];
    assign inter_7[773] = inter_6[773]^inter_6[837];
    assign inter_7[774] = inter_6[774]^inter_6[838];
    assign inter_7[775] = inter_6[775]^inter_6[839];
    assign inter_7[776] = inter_6[776]^inter_6[840];
    assign inter_7[777] = inter_6[777]^inter_6[841];
    assign inter_7[778] = inter_6[778]^inter_6[842];
    assign inter_7[779] = inter_6[779]^inter_6[843];
    assign inter_7[780] = inter_6[780]^inter_6[844];
    assign inter_7[781] = inter_6[781]^inter_6[845];
    assign inter_7[782] = inter_6[782]^inter_6[846];
    assign inter_7[783] = inter_6[783]^inter_6[847];
    assign inter_7[784] = inter_6[784]^inter_6[848];
    assign inter_7[785] = inter_6[785]^inter_6[849];
    assign inter_7[786] = inter_6[786]^inter_6[850];
    assign inter_7[787] = inter_6[787]^inter_6[851];
    assign inter_7[788] = inter_6[788]^inter_6[852];
    assign inter_7[789] = inter_6[789]^inter_6[853];
    assign inter_7[790] = inter_6[790]^inter_6[854];
    assign inter_7[791] = inter_6[791]^inter_6[855];
    assign inter_7[792] = inter_6[792]^inter_6[856];
    assign inter_7[793] = inter_6[793]^inter_6[857];
    assign inter_7[794] = inter_6[794]^inter_6[858];
    assign inter_7[795] = inter_6[795]^inter_6[859];
    assign inter_7[796] = inter_6[796]^inter_6[860];
    assign inter_7[797] = inter_6[797]^inter_6[861];
    assign inter_7[798] = inter_6[798]^inter_6[862];
    assign inter_7[799] = inter_6[799]^inter_6[863];
    assign inter_7[800] = inter_6[800]^inter_6[864];
    assign inter_7[801] = inter_6[801]^inter_6[865];
    assign inter_7[802] = inter_6[802]^inter_6[866];
    assign inter_7[803] = inter_6[803]^inter_6[867];
    assign inter_7[804] = inter_6[804]^inter_6[868];
    assign inter_7[805] = inter_6[805]^inter_6[869];
    assign inter_7[806] = inter_6[806]^inter_6[870];
    assign inter_7[807] = inter_6[807]^inter_6[871];
    assign inter_7[808] = inter_6[808]^inter_6[872];
    assign inter_7[809] = inter_6[809]^inter_6[873];
    assign inter_7[810] = inter_6[810]^inter_6[874];
    assign inter_7[811] = inter_6[811]^inter_6[875];
    assign inter_7[812] = inter_6[812]^inter_6[876];
    assign inter_7[813] = inter_6[813]^inter_6[877];
    assign inter_7[814] = inter_6[814]^inter_6[878];
    assign inter_7[815] = inter_6[815]^inter_6[879];
    assign inter_7[816] = inter_6[816]^inter_6[880];
    assign inter_7[817] = inter_6[817]^inter_6[881];
    assign inter_7[818] = inter_6[818]^inter_6[882];
    assign inter_7[819] = inter_6[819]^inter_6[883];
    assign inter_7[820] = inter_6[820]^inter_6[884];
    assign inter_7[821] = inter_6[821]^inter_6[885];
    assign inter_7[822] = inter_6[822]^inter_6[886];
    assign inter_7[823] = inter_6[823]^inter_6[887];
    assign inter_7[824] = inter_6[824]^inter_6[888];
    assign inter_7[825] = inter_6[825]^inter_6[889];
    assign inter_7[826] = inter_6[826]^inter_6[890];
    assign inter_7[827] = inter_6[827]^inter_6[891];
    assign inter_7[828] = inter_6[828]^inter_6[892];
    assign inter_7[829] = inter_6[829]^inter_6[893];
    assign inter_7[830] = inter_6[830]^inter_6[894];
    assign inter_7[831] = inter_6[831]^inter_6[895];
    assign inter_7[832] = inter_6[832];
    assign inter_7[833] = inter_6[833];
    assign inter_7[834] = inter_6[834];
    assign inter_7[835] = inter_6[835];
    assign inter_7[836] = inter_6[836];
    assign inter_7[837] = inter_6[837];
    assign inter_7[838] = inter_6[838];
    assign inter_7[839] = inter_6[839];
    assign inter_7[840] = inter_6[840];
    assign inter_7[841] = inter_6[841];
    assign inter_7[842] = inter_6[842];
    assign inter_7[843] = inter_6[843];
    assign inter_7[844] = inter_6[844];
    assign inter_7[845] = inter_6[845];
    assign inter_7[846] = inter_6[846];
    assign inter_7[847] = inter_6[847];
    assign inter_7[848] = inter_6[848];
    assign inter_7[849] = inter_6[849];
    assign inter_7[850] = inter_6[850];
    assign inter_7[851] = inter_6[851];
    assign inter_7[852] = inter_6[852];
    assign inter_7[853] = inter_6[853];
    assign inter_7[854] = inter_6[854];
    assign inter_7[855] = inter_6[855];
    assign inter_7[856] = inter_6[856];
    assign inter_7[857] = inter_6[857];
    assign inter_7[858] = inter_6[858];
    assign inter_7[859] = inter_6[859];
    assign inter_7[860] = inter_6[860];
    assign inter_7[861] = inter_6[861];
    assign inter_7[862] = inter_6[862];
    assign inter_7[863] = inter_6[863];
    assign inter_7[864] = inter_6[864];
    assign inter_7[865] = inter_6[865];
    assign inter_7[866] = inter_6[866];
    assign inter_7[867] = inter_6[867];
    assign inter_7[868] = inter_6[868];
    assign inter_7[869] = inter_6[869];
    assign inter_7[870] = inter_6[870];
    assign inter_7[871] = inter_6[871];
    assign inter_7[872] = inter_6[872];
    assign inter_7[873] = inter_6[873];
    assign inter_7[874] = inter_6[874];
    assign inter_7[875] = inter_6[875];
    assign inter_7[876] = inter_6[876];
    assign inter_7[877] = inter_6[877];
    assign inter_7[878] = inter_6[878];
    assign inter_7[879] = inter_6[879];
    assign inter_7[880] = inter_6[880];
    assign inter_7[881] = inter_6[881];
    assign inter_7[882] = inter_6[882];
    assign inter_7[883] = inter_6[883];
    assign inter_7[884] = inter_6[884];
    assign inter_7[885] = inter_6[885];
    assign inter_7[886] = inter_6[886];
    assign inter_7[887] = inter_6[887];
    assign inter_7[888] = inter_6[888];
    assign inter_7[889] = inter_6[889];
    assign inter_7[890] = inter_6[890];
    assign inter_7[891] = inter_6[891];
    assign inter_7[892] = inter_6[892];
    assign inter_7[893] = inter_6[893];
    assign inter_7[894] = inter_6[894];
    assign inter_7[895] = inter_6[895];
    assign inter_7[896] = inter_6[896]^inter_6[960];
    assign inter_7[897] = inter_6[897]^inter_6[961];
    assign inter_7[898] = inter_6[898]^inter_6[962];
    assign inter_7[899] = inter_6[899]^inter_6[963];
    assign inter_7[900] = inter_6[900]^inter_6[964];
    assign inter_7[901] = inter_6[901]^inter_6[965];
    assign inter_7[902] = inter_6[902]^inter_6[966];
    assign inter_7[903] = inter_6[903]^inter_6[967];
    assign inter_7[904] = inter_6[904]^inter_6[968];
    assign inter_7[905] = inter_6[905]^inter_6[969];
    assign inter_7[906] = inter_6[906]^inter_6[970];
    assign inter_7[907] = inter_6[907]^inter_6[971];
    assign inter_7[908] = inter_6[908]^inter_6[972];
    assign inter_7[909] = inter_6[909]^inter_6[973];
    assign inter_7[910] = inter_6[910]^inter_6[974];
    assign inter_7[911] = inter_6[911]^inter_6[975];
    assign inter_7[912] = inter_6[912]^inter_6[976];
    assign inter_7[913] = inter_6[913]^inter_6[977];
    assign inter_7[914] = inter_6[914]^inter_6[978];
    assign inter_7[915] = inter_6[915]^inter_6[979];
    assign inter_7[916] = inter_6[916]^inter_6[980];
    assign inter_7[917] = inter_6[917]^inter_6[981];
    assign inter_7[918] = inter_6[918]^inter_6[982];
    assign inter_7[919] = inter_6[919]^inter_6[983];
    assign inter_7[920] = inter_6[920]^inter_6[984];
    assign inter_7[921] = inter_6[921]^inter_6[985];
    assign inter_7[922] = inter_6[922]^inter_6[986];
    assign inter_7[923] = inter_6[923]^inter_6[987];
    assign inter_7[924] = inter_6[924]^inter_6[988];
    assign inter_7[925] = inter_6[925]^inter_6[989];
    assign inter_7[926] = inter_6[926]^inter_6[990];
    assign inter_7[927] = inter_6[927]^inter_6[991];
    assign inter_7[928] = inter_6[928]^inter_6[992];
    assign inter_7[929] = inter_6[929]^inter_6[993];
    assign inter_7[930] = inter_6[930]^inter_6[994];
    assign inter_7[931] = inter_6[931]^inter_6[995];
    assign inter_7[932] = inter_6[932]^inter_6[996];
    assign inter_7[933] = inter_6[933]^inter_6[997];
    assign inter_7[934] = inter_6[934]^inter_6[998];
    assign inter_7[935] = inter_6[935]^inter_6[999];
    assign inter_7[936] = inter_6[936]^inter_6[1000];
    assign inter_7[937] = inter_6[937]^inter_6[1001];
    assign inter_7[938] = inter_6[938]^inter_6[1002];
    assign inter_7[939] = inter_6[939]^inter_6[1003];
    assign inter_7[940] = inter_6[940]^inter_6[1004];
    assign inter_7[941] = inter_6[941]^inter_6[1005];
    assign inter_7[942] = inter_6[942]^inter_6[1006];
    assign inter_7[943] = inter_6[943]^inter_6[1007];
    assign inter_7[944] = inter_6[944]^inter_6[1008];
    assign inter_7[945] = inter_6[945]^inter_6[1009];
    assign inter_7[946] = inter_6[946]^inter_6[1010];
    assign inter_7[947] = inter_6[947]^inter_6[1011];
    assign inter_7[948] = inter_6[948]^inter_6[1012];
    assign inter_7[949] = inter_6[949]^inter_6[1013];
    assign inter_7[950] = inter_6[950]^inter_6[1014];
    assign inter_7[951] = inter_6[951]^inter_6[1015];
    assign inter_7[952] = inter_6[952]^inter_6[1016];
    assign inter_7[953] = inter_6[953]^inter_6[1017];
    assign inter_7[954] = inter_6[954]^inter_6[1018];
    assign inter_7[955] = inter_6[955]^inter_6[1019];
    assign inter_7[956] = inter_6[956]^inter_6[1020];
    assign inter_7[957] = inter_6[957]^inter_6[1021];
    assign inter_7[958] = inter_6[958]^inter_6[1022];
    assign inter_7[959] = inter_6[959]^inter_6[1023];
    assign inter_7[960] = inter_6[960];
    assign inter_7[961] = inter_6[961];
    assign inter_7[962] = inter_6[962];
    assign inter_7[963] = inter_6[963];
    assign inter_7[964] = inter_6[964];
    assign inter_7[965] = inter_6[965];
    assign inter_7[966] = inter_6[966];
    assign inter_7[967] = inter_6[967];
    assign inter_7[968] = inter_6[968];
    assign inter_7[969] = inter_6[969];
    assign inter_7[970] = inter_6[970];
    assign inter_7[971] = inter_6[971];
    assign inter_7[972] = inter_6[972];
    assign inter_7[973] = inter_6[973];
    assign inter_7[974] = inter_6[974];
    assign inter_7[975] = inter_6[975];
    assign inter_7[976] = inter_6[976];
    assign inter_7[977] = inter_6[977];
    assign inter_7[978] = inter_6[978];
    assign inter_7[979] = inter_6[979];
    assign inter_7[980] = inter_6[980];
    assign inter_7[981] = inter_6[981];
    assign inter_7[982] = inter_6[982];
    assign inter_7[983] = inter_6[983];
    assign inter_7[984] = inter_6[984];
    assign inter_7[985] = inter_6[985];
    assign inter_7[986] = inter_6[986];
    assign inter_7[987] = inter_6[987];
    assign inter_7[988] = inter_6[988];
    assign inter_7[989] = inter_6[989];
    assign inter_7[990] = inter_6[990];
    assign inter_7[991] = inter_6[991];
    assign inter_7[992] = inter_6[992];
    assign inter_7[993] = inter_6[993];
    assign inter_7[994] = inter_6[994];
    assign inter_7[995] = inter_6[995];
    assign inter_7[996] = inter_6[996];
    assign inter_7[997] = inter_6[997];
    assign inter_7[998] = inter_6[998];
    assign inter_7[999] = inter_6[999];
    assign inter_7[1000] = inter_6[1000];
    assign inter_7[1001] = inter_6[1001];
    assign inter_7[1002] = inter_6[1002];
    assign inter_7[1003] = inter_6[1003];
    assign inter_7[1004] = inter_6[1004];
    assign inter_7[1005] = inter_6[1005];
    assign inter_7[1006] = inter_6[1006];
    assign inter_7[1007] = inter_6[1007];
    assign inter_7[1008] = inter_6[1008];
    assign inter_7[1009] = inter_6[1009];
    assign inter_7[1010] = inter_6[1010];
    assign inter_7[1011] = inter_6[1011];
    assign inter_7[1012] = inter_6[1012];
    assign inter_7[1013] = inter_6[1013];
    assign inter_7[1014] = inter_6[1014];
    assign inter_7[1015] = inter_6[1015];
    assign inter_7[1016] = inter_6[1016];
    assign inter_7[1017] = inter_6[1017];
    assign inter_7[1018] = inter_6[1018];
    assign inter_7[1019] = inter_6[1019];
    assign inter_7[1020] = inter_6[1020];
    assign inter_7[1021] = inter_6[1021];
    assign inter_7[1022] = inter_6[1022];
    assign inter_7[1023] = inter_6[1023];
    /***************************/
    assign inter_8[0] = inter_7[0]^inter_7[128];
    assign inter_8[1] = inter_7[1]^inter_7[129];
    assign inter_8[2] = inter_7[2]^inter_7[130];
    assign inter_8[3] = inter_7[3]^inter_7[131];
    assign inter_8[4] = inter_7[4]^inter_7[132];
    assign inter_8[5] = inter_7[5]^inter_7[133];
    assign inter_8[6] = inter_7[6]^inter_7[134];
    assign inter_8[7] = inter_7[7]^inter_7[135];
    assign inter_8[8] = inter_7[8]^inter_7[136];
    assign inter_8[9] = inter_7[9]^inter_7[137];
    assign inter_8[10] = inter_7[10]^inter_7[138];
    assign inter_8[11] = inter_7[11]^inter_7[139];
    assign inter_8[12] = inter_7[12]^inter_7[140];
    assign inter_8[13] = inter_7[13]^inter_7[141];
    assign inter_8[14] = inter_7[14]^inter_7[142];
    assign inter_8[15] = inter_7[15]^inter_7[143];
    assign inter_8[16] = inter_7[16]^inter_7[144];
    assign inter_8[17] = inter_7[17]^inter_7[145];
    assign inter_8[18] = inter_7[18]^inter_7[146];
    assign inter_8[19] = inter_7[19]^inter_7[147];
    assign inter_8[20] = inter_7[20]^inter_7[148];
    assign inter_8[21] = inter_7[21]^inter_7[149];
    assign inter_8[22] = inter_7[22]^inter_7[150];
    assign inter_8[23] = inter_7[23]^inter_7[151];
    assign inter_8[24] = inter_7[24]^inter_7[152];
    assign inter_8[25] = inter_7[25]^inter_7[153];
    assign inter_8[26] = inter_7[26]^inter_7[154];
    assign inter_8[27] = inter_7[27]^inter_7[155];
    assign inter_8[28] = inter_7[28]^inter_7[156];
    assign inter_8[29] = inter_7[29]^inter_7[157];
    assign inter_8[30] = inter_7[30]^inter_7[158];
    assign inter_8[31] = inter_7[31]^inter_7[159];
    assign inter_8[32] = inter_7[32]^inter_7[160];
    assign inter_8[33] = inter_7[33]^inter_7[161];
    assign inter_8[34] = inter_7[34]^inter_7[162];
    assign inter_8[35] = inter_7[35]^inter_7[163];
    assign inter_8[36] = inter_7[36]^inter_7[164];
    assign inter_8[37] = inter_7[37]^inter_7[165];
    assign inter_8[38] = inter_7[38]^inter_7[166];
    assign inter_8[39] = inter_7[39]^inter_7[167];
    assign inter_8[40] = inter_7[40]^inter_7[168];
    assign inter_8[41] = inter_7[41]^inter_7[169];
    assign inter_8[42] = inter_7[42]^inter_7[170];
    assign inter_8[43] = inter_7[43]^inter_7[171];
    assign inter_8[44] = inter_7[44]^inter_7[172];
    assign inter_8[45] = inter_7[45]^inter_7[173];
    assign inter_8[46] = inter_7[46]^inter_7[174];
    assign inter_8[47] = inter_7[47]^inter_7[175];
    assign inter_8[48] = inter_7[48]^inter_7[176];
    assign inter_8[49] = inter_7[49]^inter_7[177];
    assign inter_8[50] = inter_7[50]^inter_7[178];
    assign inter_8[51] = inter_7[51]^inter_7[179];
    assign inter_8[52] = inter_7[52]^inter_7[180];
    assign inter_8[53] = inter_7[53]^inter_7[181];
    assign inter_8[54] = inter_7[54]^inter_7[182];
    assign inter_8[55] = inter_7[55]^inter_7[183];
    assign inter_8[56] = inter_7[56]^inter_7[184];
    assign inter_8[57] = inter_7[57]^inter_7[185];
    assign inter_8[58] = inter_7[58]^inter_7[186];
    assign inter_8[59] = inter_7[59]^inter_7[187];
    assign inter_8[60] = inter_7[60]^inter_7[188];
    assign inter_8[61] = inter_7[61]^inter_7[189];
    assign inter_8[62] = inter_7[62]^inter_7[190];
    assign inter_8[63] = inter_7[63]^inter_7[191];
    assign inter_8[64] = inter_7[64]^inter_7[192];
    assign inter_8[65] = inter_7[65]^inter_7[193];
    assign inter_8[66] = inter_7[66]^inter_7[194];
    assign inter_8[67] = inter_7[67]^inter_7[195];
    assign inter_8[68] = inter_7[68]^inter_7[196];
    assign inter_8[69] = inter_7[69]^inter_7[197];
    assign inter_8[70] = inter_7[70]^inter_7[198];
    assign inter_8[71] = inter_7[71]^inter_7[199];
    assign inter_8[72] = inter_7[72]^inter_7[200];
    assign inter_8[73] = inter_7[73]^inter_7[201];
    assign inter_8[74] = inter_7[74]^inter_7[202];
    assign inter_8[75] = inter_7[75]^inter_7[203];
    assign inter_8[76] = inter_7[76]^inter_7[204];
    assign inter_8[77] = inter_7[77]^inter_7[205];
    assign inter_8[78] = inter_7[78]^inter_7[206];
    assign inter_8[79] = inter_7[79]^inter_7[207];
    assign inter_8[80] = inter_7[80]^inter_7[208];
    assign inter_8[81] = inter_7[81]^inter_7[209];
    assign inter_8[82] = inter_7[82]^inter_7[210];
    assign inter_8[83] = inter_7[83]^inter_7[211];
    assign inter_8[84] = inter_7[84]^inter_7[212];
    assign inter_8[85] = inter_7[85]^inter_7[213];
    assign inter_8[86] = inter_7[86]^inter_7[214];
    assign inter_8[87] = inter_7[87]^inter_7[215];
    assign inter_8[88] = inter_7[88]^inter_7[216];
    assign inter_8[89] = inter_7[89]^inter_7[217];
    assign inter_8[90] = inter_7[90]^inter_7[218];
    assign inter_8[91] = inter_7[91]^inter_7[219];
    assign inter_8[92] = inter_7[92]^inter_7[220];
    assign inter_8[93] = inter_7[93]^inter_7[221];
    assign inter_8[94] = inter_7[94]^inter_7[222];
    assign inter_8[95] = inter_7[95]^inter_7[223];
    assign inter_8[96] = inter_7[96]^inter_7[224];
    assign inter_8[97] = inter_7[97]^inter_7[225];
    assign inter_8[98] = inter_7[98]^inter_7[226];
    assign inter_8[99] = inter_7[99]^inter_7[227];
    assign inter_8[100] = inter_7[100]^inter_7[228];
    assign inter_8[101] = inter_7[101]^inter_7[229];
    assign inter_8[102] = inter_7[102]^inter_7[230];
    assign inter_8[103] = inter_7[103]^inter_7[231];
    assign inter_8[104] = inter_7[104]^inter_7[232];
    assign inter_8[105] = inter_7[105]^inter_7[233];
    assign inter_8[106] = inter_7[106]^inter_7[234];
    assign inter_8[107] = inter_7[107]^inter_7[235];
    assign inter_8[108] = inter_7[108]^inter_7[236];
    assign inter_8[109] = inter_7[109]^inter_7[237];
    assign inter_8[110] = inter_7[110]^inter_7[238];
    assign inter_8[111] = inter_7[111]^inter_7[239];
    assign inter_8[112] = inter_7[112]^inter_7[240];
    assign inter_8[113] = inter_7[113]^inter_7[241];
    assign inter_8[114] = inter_7[114]^inter_7[242];
    assign inter_8[115] = inter_7[115]^inter_7[243];
    assign inter_8[116] = inter_7[116]^inter_7[244];
    assign inter_8[117] = inter_7[117]^inter_7[245];
    assign inter_8[118] = inter_7[118]^inter_7[246];
    assign inter_8[119] = inter_7[119]^inter_7[247];
    assign inter_8[120] = inter_7[120]^inter_7[248];
    assign inter_8[121] = inter_7[121]^inter_7[249];
    assign inter_8[122] = inter_7[122]^inter_7[250];
    assign inter_8[123] = inter_7[123]^inter_7[251];
    assign inter_8[124] = inter_7[124]^inter_7[252];
    assign inter_8[125] = inter_7[125]^inter_7[253];
    assign inter_8[126] = inter_7[126]^inter_7[254];
    assign inter_8[127] = inter_7[127]^inter_7[255];
    assign inter_8[128] = inter_7[128];
    assign inter_8[129] = inter_7[129];
    assign inter_8[130] = inter_7[130];
    assign inter_8[131] = inter_7[131];
    assign inter_8[132] = inter_7[132];
    assign inter_8[133] = inter_7[133];
    assign inter_8[134] = inter_7[134];
    assign inter_8[135] = inter_7[135];
    assign inter_8[136] = inter_7[136];
    assign inter_8[137] = inter_7[137];
    assign inter_8[138] = inter_7[138];
    assign inter_8[139] = inter_7[139];
    assign inter_8[140] = inter_7[140];
    assign inter_8[141] = inter_7[141];
    assign inter_8[142] = inter_7[142];
    assign inter_8[143] = inter_7[143];
    assign inter_8[144] = inter_7[144];
    assign inter_8[145] = inter_7[145];
    assign inter_8[146] = inter_7[146];
    assign inter_8[147] = inter_7[147];
    assign inter_8[148] = inter_7[148];
    assign inter_8[149] = inter_7[149];
    assign inter_8[150] = inter_7[150];
    assign inter_8[151] = inter_7[151];
    assign inter_8[152] = inter_7[152];
    assign inter_8[153] = inter_7[153];
    assign inter_8[154] = inter_7[154];
    assign inter_8[155] = inter_7[155];
    assign inter_8[156] = inter_7[156];
    assign inter_8[157] = inter_7[157];
    assign inter_8[158] = inter_7[158];
    assign inter_8[159] = inter_7[159];
    assign inter_8[160] = inter_7[160];
    assign inter_8[161] = inter_7[161];
    assign inter_8[162] = inter_7[162];
    assign inter_8[163] = inter_7[163];
    assign inter_8[164] = inter_7[164];
    assign inter_8[165] = inter_7[165];
    assign inter_8[166] = inter_7[166];
    assign inter_8[167] = inter_7[167];
    assign inter_8[168] = inter_7[168];
    assign inter_8[169] = inter_7[169];
    assign inter_8[170] = inter_7[170];
    assign inter_8[171] = inter_7[171];
    assign inter_8[172] = inter_7[172];
    assign inter_8[173] = inter_7[173];
    assign inter_8[174] = inter_7[174];
    assign inter_8[175] = inter_7[175];
    assign inter_8[176] = inter_7[176];
    assign inter_8[177] = inter_7[177];
    assign inter_8[178] = inter_7[178];
    assign inter_8[179] = inter_7[179];
    assign inter_8[180] = inter_7[180];
    assign inter_8[181] = inter_7[181];
    assign inter_8[182] = inter_7[182];
    assign inter_8[183] = inter_7[183];
    assign inter_8[184] = inter_7[184];
    assign inter_8[185] = inter_7[185];
    assign inter_8[186] = inter_7[186];
    assign inter_8[187] = inter_7[187];
    assign inter_8[188] = inter_7[188];
    assign inter_8[189] = inter_7[189];
    assign inter_8[190] = inter_7[190];
    assign inter_8[191] = inter_7[191];
    assign inter_8[192] = inter_7[192];
    assign inter_8[193] = inter_7[193];
    assign inter_8[194] = inter_7[194];
    assign inter_8[195] = inter_7[195];
    assign inter_8[196] = inter_7[196];
    assign inter_8[197] = inter_7[197];
    assign inter_8[198] = inter_7[198];
    assign inter_8[199] = inter_7[199];
    assign inter_8[200] = inter_7[200];
    assign inter_8[201] = inter_7[201];
    assign inter_8[202] = inter_7[202];
    assign inter_8[203] = inter_7[203];
    assign inter_8[204] = inter_7[204];
    assign inter_8[205] = inter_7[205];
    assign inter_8[206] = inter_7[206];
    assign inter_8[207] = inter_7[207];
    assign inter_8[208] = inter_7[208];
    assign inter_8[209] = inter_7[209];
    assign inter_8[210] = inter_7[210];
    assign inter_8[211] = inter_7[211];
    assign inter_8[212] = inter_7[212];
    assign inter_8[213] = inter_7[213];
    assign inter_8[214] = inter_7[214];
    assign inter_8[215] = inter_7[215];
    assign inter_8[216] = inter_7[216];
    assign inter_8[217] = inter_7[217];
    assign inter_8[218] = inter_7[218];
    assign inter_8[219] = inter_7[219];
    assign inter_8[220] = inter_7[220];
    assign inter_8[221] = inter_7[221];
    assign inter_8[222] = inter_7[222];
    assign inter_8[223] = inter_7[223];
    assign inter_8[224] = inter_7[224];
    assign inter_8[225] = inter_7[225];
    assign inter_8[226] = inter_7[226];
    assign inter_8[227] = inter_7[227];
    assign inter_8[228] = inter_7[228];
    assign inter_8[229] = inter_7[229];
    assign inter_8[230] = inter_7[230];
    assign inter_8[231] = inter_7[231];
    assign inter_8[232] = inter_7[232];
    assign inter_8[233] = inter_7[233];
    assign inter_8[234] = inter_7[234];
    assign inter_8[235] = inter_7[235];
    assign inter_8[236] = inter_7[236];
    assign inter_8[237] = inter_7[237];
    assign inter_8[238] = inter_7[238];
    assign inter_8[239] = inter_7[239];
    assign inter_8[240] = inter_7[240];
    assign inter_8[241] = inter_7[241];
    assign inter_8[242] = inter_7[242];
    assign inter_8[243] = inter_7[243];
    assign inter_8[244] = inter_7[244];
    assign inter_8[245] = inter_7[245];
    assign inter_8[246] = inter_7[246];
    assign inter_8[247] = inter_7[247];
    assign inter_8[248] = inter_7[248];
    assign inter_8[249] = inter_7[249];
    assign inter_8[250] = inter_7[250];
    assign inter_8[251] = inter_7[251];
    assign inter_8[252] = inter_7[252];
    assign inter_8[253] = inter_7[253];
    assign inter_8[254] = inter_7[254];
    assign inter_8[255] = inter_7[255];
    assign inter_8[256] = inter_7[256]^inter_7[384];
    assign inter_8[257] = inter_7[257]^inter_7[385];
    assign inter_8[258] = inter_7[258]^inter_7[386];
    assign inter_8[259] = inter_7[259]^inter_7[387];
    assign inter_8[260] = inter_7[260]^inter_7[388];
    assign inter_8[261] = inter_7[261]^inter_7[389];
    assign inter_8[262] = inter_7[262]^inter_7[390];
    assign inter_8[263] = inter_7[263]^inter_7[391];
    assign inter_8[264] = inter_7[264]^inter_7[392];
    assign inter_8[265] = inter_7[265]^inter_7[393];
    assign inter_8[266] = inter_7[266]^inter_7[394];
    assign inter_8[267] = inter_7[267]^inter_7[395];
    assign inter_8[268] = inter_7[268]^inter_7[396];
    assign inter_8[269] = inter_7[269]^inter_7[397];
    assign inter_8[270] = inter_7[270]^inter_7[398];
    assign inter_8[271] = inter_7[271]^inter_7[399];
    assign inter_8[272] = inter_7[272]^inter_7[400];
    assign inter_8[273] = inter_7[273]^inter_7[401];
    assign inter_8[274] = inter_7[274]^inter_7[402];
    assign inter_8[275] = inter_7[275]^inter_7[403];
    assign inter_8[276] = inter_7[276]^inter_7[404];
    assign inter_8[277] = inter_7[277]^inter_7[405];
    assign inter_8[278] = inter_7[278]^inter_7[406];
    assign inter_8[279] = inter_7[279]^inter_7[407];
    assign inter_8[280] = inter_7[280]^inter_7[408];
    assign inter_8[281] = inter_7[281]^inter_7[409];
    assign inter_8[282] = inter_7[282]^inter_7[410];
    assign inter_8[283] = inter_7[283]^inter_7[411];
    assign inter_8[284] = inter_7[284]^inter_7[412];
    assign inter_8[285] = inter_7[285]^inter_7[413];
    assign inter_8[286] = inter_7[286]^inter_7[414];
    assign inter_8[287] = inter_7[287]^inter_7[415];
    assign inter_8[288] = inter_7[288]^inter_7[416];
    assign inter_8[289] = inter_7[289]^inter_7[417];
    assign inter_8[290] = inter_7[290]^inter_7[418];
    assign inter_8[291] = inter_7[291]^inter_7[419];
    assign inter_8[292] = inter_7[292]^inter_7[420];
    assign inter_8[293] = inter_7[293]^inter_7[421];
    assign inter_8[294] = inter_7[294]^inter_7[422];
    assign inter_8[295] = inter_7[295]^inter_7[423];
    assign inter_8[296] = inter_7[296]^inter_7[424];
    assign inter_8[297] = inter_7[297]^inter_7[425];
    assign inter_8[298] = inter_7[298]^inter_7[426];
    assign inter_8[299] = inter_7[299]^inter_7[427];
    assign inter_8[300] = inter_7[300]^inter_7[428];
    assign inter_8[301] = inter_7[301]^inter_7[429];
    assign inter_8[302] = inter_7[302]^inter_7[430];
    assign inter_8[303] = inter_7[303]^inter_7[431];
    assign inter_8[304] = inter_7[304]^inter_7[432];
    assign inter_8[305] = inter_7[305]^inter_7[433];
    assign inter_8[306] = inter_7[306]^inter_7[434];
    assign inter_8[307] = inter_7[307]^inter_7[435];
    assign inter_8[308] = inter_7[308]^inter_7[436];
    assign inter_8[309] = inter_7[309]^inter_7[437];
    assign inter_8[310] = inter_7[310]^inter_7[438];
    assign inter_8[311] = inter_7[311]^inter_7[439];
    assign inter_8[312] = inter_7[312]^inter_7[440];
    assign inter_8[313] = inter_7[313]^inter_7[441];
    assign inter_8[314] = inter_7[314]^inter_7[442];
    assign inter_8[315] = inter_7[315]^inter_7[443];
    assign inter_8[316] = inter_7[316]^inter_7[444];
    assign inter_8[317] = inter_7[317]^inter_7[445];
    assign inter_8[318] = inter_7[318]^inter_7[446];
    assign inter_8[319] = inter_7[319]^inter_7[447];
    assign inter_8[320] = inter_7[320]^inter_7[448];
    assign inter_8[321] = inter_7[321]^inter_7[449];
    assign inter_8[322] = inter_7[322]^inter_7[450];
    assign inter_8[323] = inter_7[323]^inter_7[451];
    assign inter_8[324] = inter_7[324]^inter_7[452];
    assign inter_8[325] = inter_7[325]^inter_7[453];
    assign inter_8[326] = inter_7[326]^inter_7[454];
    assign inter_8[327] = inter_7[327]^inter_7[455];
    assign inter_8[328] = inter_7[328]^inter_7[456];
    assign inter_8[329] = inter_7[329]^inter_7[457];
    assign inter_8[330] = inter_7[330]^inter_7[458];
    assign inter_8[331] = inter_7[331]^inter_7[459];
    assign inter_8[332] = inter_7[332]^inter_7[460];
    assign inter_8[333] = inter_7[333]^inter_7[461];
    assign inter_8[334] = inter_7[334]^inter_7[462];
    assign inter_8[335] = inter_7[335]^inter_7[463];
    assign inter_8[336] = inter_7[336]^inter_7[464];
    assign inter_8[337] = inter_7[337]^inter_7[465];
    assign inter_8[338] = inter_7[338]^inter_7[466];
    assign inter_8[339] = inter_7[339]^inter_7[467];
    assign inter_8[340] = inter_7[340]^inter_7[468];
    assign inter_8[341] = inter_7[341]^inter_7[469];
    assign inter_8[342] = inter_7[342]^inter_7[470];
    assign inter_8[343] = inter_7[343]^inter_7[471];
    assign inter_8[344] = inter_7[344]^inter_7[472];
    assign inter_8[345] = inter_7[345]^inter_7[473];
    assign inter_8[346] = inter_7[346]^inter_7[474];
    assign inter_8[347] = inter_7[347]^inter_7[475];
    assign inter_8[348] = inter_7[348]^inter_7[476];
    assign inter_8[349] = inter_7[349]^inter_7[477];
    assign inter_8[350] = inter_7[350]^inter_7[478];
    assign inter_8[351] = inter_7[351]^inter_7[479];
    assign inter_8[352] = inter_7[352]^inter_7[480];
    assign inter_8[353] = inter_7[353]^inter_7[481];
    assign inter_8[354] = inter_7[354]^inter_7[482];
    assign inter_8[355] = inter_7[355]^inter_7[483];
    assign inter_8[356] = inter_7[356]^inter_7[484];
    assign inter_8[357] = inter_7[357]^inter_7[485];
    assign inter_8[358] = inter_7[358]^inter_7[486];
    assign inter_8[359] = inter_7[359]^inter_7[487];
    assign inter_8[360] = inter_7[360]^inter_7[488];
    assign inter_8[361] = inter_7[361]^inter_7[489];
    assign inter_8[362] = inter_7[362]^inter_7[490];
    assign inter_8[363] = inter_7[363]^inter_7[491];
    assign inter_8[364] = inter_7[364]^inter_7[492];
    assign inter_8[365] = inter_7[365]^inter_7[493];
    assign inter_8[366] = inter_7[366]^inter_7[494];
    assign inter_8[367] = inter_7[367]^inter_7[495];
    assign inter_8[368] = inter_7[368]^inter_7[496];
    assign inter_8[369] = inter_7[369]^inter_7[497];
    assign inter_8[370] = inter_7[370]^inter_7[498];
    assign inter_8[371] = inter_7[371]^inter_7[499];
    assign inter_8[372] = inter_7[372]^inter_7[500];
    assign inter_8[373] = inter_7[373]^inter_7[501];
    assign inter_8[374] = inter_7[374]^inter_7[502];
    assign inter_8[375] = inter_7[375]^inter_7[503];
    assign inter_8[376] = inter_7[376]^inter_7[504];
    assign inter_8[377] = inter_7[377]^inter_7[505];
    assign inter_8[378] = inter_7[378]^inter_7[506];
    assign inter_8[379] = inter_7[379]^inter_7[507];
    assign inter_8[380] = inter_7[380]^inter_7[508];
    assign inter_8[381] = inter_7[381]^inter_7[509];
    assign inter_8[382] = inter_7[382]^inter_7[510];
    assign inter_8[383] = inter_7[383]^inter_7[511];
    assign inter_8[384] = inter_7[384];
    assign inter_8[385] = inter_7[385];
    assign inter_8[386] = inter_7[386];
    assign inter_8[387] = inter_7[387];
    assign inter_8[388] = inter_7[388];
    assign inter_8[389] = inter_7[389];
    assign inter_8[390] = inter_7[390];
    assign inter_8[391] = inter_7[391];
    assign inter_8[392] = inter_7[392];
    assign inter_8[393] = inter_7[393];
    assign inter_8[394] = inter_7[394];
    assign inter_8[395] = inter_7[395];
    assign inter_8[396] = inter_7[396];
    assign inter_8[397] = inter_7[397];
    assign inter_8[398] = inter_7[398];
    assign inter_8[399] = inter_7[399];
    assign inter_8[400] = inter_7[400];
    assign inter_8[401] = inter_7[401];
    assign inter_8[402] = inter_7[402];
    assign inter_8[403] = inter_7[403];
    assign inter_8[404] = inter_7[404];
    assign inter_8[405] = inter_7[405];
    assign inter_8[406] = inter_7[406];
    assign inter_8[407] = inter_7[407];
    assign inter_8[408] = inter_7[408];
    assign inter_8[409] = inter_7[409];
    assign inter_8[410] = inter_7[410];
    assign inter_8[411] = inter_7[411];
    assign inter_8[412] = inter_7[412];
    assign inter_8[413] = inter_7[413];
    assign inter_8[414] = inter_7[414];
    assign inter_8[415] = inter_7[415];
    assign inter_8[416] = inter_7[416];
    assign inter_8[417] = inter_7[417];
    assign inter_8[418] = inter_7[418];
    assign inter_8[419] = inter_7[419];
    assign inter_8[420] = inter_7[420];
    assign inter_8[421] = inter_7[421];
    assign inter_8[422] = inter_7[422];
    assign inter_8[423] = inter_7[423];
    assign inter_8[424] = inter_7[424];
    assign inter_8[425] = inter_7[425];
    assign inter_8[426] = inter_7[426];
    assign inter_8[427] = inter_7[427];
    assign inter_8[428] = inter_7[428];
    assign inter_8[429] = inter_7[429];
    assign inter_8[430] = inter_7[430];
    assign inter_8[431] = inter_7[431];
    assign inter_8[432] = inter_7[432];
    assign inter_8[433] = inter_7[433];
    assign inter_8[434] = inter_7[434];
    assign inter_8[435] = inter_7[435];
    assign inter_8[436] = inter_7[436];
    assign inter_8[437] = inter_7[437];
    assign inter_8[438] = inter_7[438];
    assign inter_8[439] = inter_7[439];
    assign inter_8[440] = inter_7[440];
    assign inter_8[441] = inter_7[441];
    assign inter_8[442] = inter_7[442];
    assign inter_8[443] = inter_7[443];
    assign inter_8[444] = inter_7[444];
    assign inter_8[445] = inter_7[445];
    assign inter_8[446] = inter_7[446];
    assign inter_8[447] = inter_7[447];
    assign inter_8[448] = inter_7[448];
    assign inter_8[449] = inter_7[449];
    assign inter_8[450] = inter_7[450];
    assign inter_8[451] = inter_7[451];
    assign inter_8[452] = inter_7[452];
    assign inter_8[453] = inter_7[453];
    assign inter_8[454] = inter_7[454];
    assign inter_8[455] = inter_7[455];
    assign inter_8[456] = inter_7[456];
    assign inter_8[457] = inter_7[457];
    assign inter_8[458] = inter_7[458];
    assign inter_8[459] = inter_7[459];
    assign inter_8[460] = inter_7[460];
    assign inter_8[461] = inter_7[461];
    assign inter_8[462] = inter_7[462];
    assign inter_8[463] = inter_7[463];
    assign inter_8[464] = inter_7[464];
    assign inter_8[465] = inter_7[465];
    assign inter_8[466] = inter_7[466];
    assign inter_8[467] = inter_7[467];
    assign inter_8[468] = inter_7[468];
    assign inter_8[469] = inter_7[469];
    assign inter_8[470] = inter_7[470];
    assign inter_8[471] = inter_7[471];
    assign inter_8[472] = inter_7[472];
    assign inter_8[473] = inter_7[473];
    assign inter_8[474] = inter_7[474];
    assign inter_8[475] = inter_7[475];
    assign inter_8[476] = inter_7[476];
    assign inter_8[477] = inter_7[477];
    assign inter_8[478] = inter_7[478];
    assign inter_8[479] = inter_7[479];
    assign inter_8[480] = inter_7[480];
    assign inter_8[481] = inter_7[481];
    assign inter_8[482] = inter_7[482];
    assign inter_8[483] = inter_7[483];
    assign inter_8[484] = inter_7[484];
    assign inter_8[485] = inter_7[485];
    assign inter_8[486] = inter_7[486];
    assign inter_8[487] = inter_7[487];
    assign inter_8[488] = inter_7[488];
    assign inter_8[489] = inter_7[489];
    assign inter_8[490] = inter_7[490];
    assign inter_8[491] = inter_7[491];
    assign inter_8[492] = inter_7[492];
    assign inter_8[493] = inter_7[493];
    assign inter_8[494] = inter_7[494];
    assign inter_8[495] = inter_7[495];
    assign inter_8[496] = inter_7[496];
    assign inter_8[497] = inter_7[497];
    assign inter_8[498] = inter_7[498];
    assign inter_8[499] = inter_7[499];
    assign inter_8[500] = inter_7[500];
    assign inter_8[501] = inter_7[501];
    assign inter_8[502] = inter_7[502];
    assign inter_8[503] = inter_7[503];
    assign inter_8[504] = inter_7[504];
    assign inter_8[505] = inter_7[505];
    assign inter_8[506] = inter_7[506];
    assign inter_8[507] = inter_7[507];
    assign inter_8[508] = inter_7[508];
    assign inter_8[509] = inter_7[509];
    assign inter_8[510] = inter_7[510];
    assign inter_8[511] = inter_7[511];
    assign inter_8[512] = inter_7[512]^inter_7[640];
    assign inter_8[513] = inter_7[513]^inter_7[641];
    assign inter_8[514] = inter_7[514]^inter_7[642];
    assign inter_8[515] = inter_7[515]^inter_7[643];
    assign inter_8[516] = inter_7[516]^inter_7[644];
    assign inter_8[517] = inter_7[517]^inter_7[645];
    assign inter_8[518] = inter_7[518]^inter_7[646];
    assign inter_8[519] = inter_7[519]^inter_7[647];
    assign inter_8[520] = inter_7[520]^inter_7[648];
    assign inter_8[521] = inter_7[521]^inter_7[649];
    assign inter_8[522] = inter_7[522]^inter_7[650];
    assign inter_8[523] = inter_7[523]^inter_7[651];
    assign inter_8[524] = inter_7[524]^inter_7[652];
    assign inter_8[525] = inter_7[525]^inter_7[653];
    assign inter_8[526] = inter_7[526]^inter_7[654];
    assign inter_8[527] = inter_7[527]^inter_7[655];
    assign inter_8[528] = inter_7[528]^inter_7[656];
    assign inter_8[529] = inter_7[529]^inter_7[657];
    assign inter_8[530] = inter_7[530]^inter_7[658];
    assign inter_8[531] = inter_7[531]^inter_7[659];
    assign inter_8[532] = inter_7[532]^inter_7[660];
    assign inter_8[533] = inter_7[533]^inter_7[661];
    assign inter_8[534] = inter_7[534]^inter_7[662];
    assign inter_8[535] = inter_7[535]^inter_7[663];
    assign inter_8[536] = inter_7[536]^inter_7[664];
    assign inter_8[537] = inter_7[537]^inter_7[665];
    assign inter_8[538] = inter_7[538]^inter_7[666];
    assign inter_8[539] = inter_7[539]^inter_7[667];
    assign inter_8[540] = inter_7[540]^inter_7[668];
    assign inter_8[541] = inter_7[541]^inter_7[669];
    assign inter_8[542] = inter_7[542]^inter_7[670];
    assign inter_8[543] = inter_7[543]^inter_7[671];
    assign inter_8[544] = inter_7[544]^inter_7[672];
    assign inter_8[545] = inter_7[545]^inter_7[673];
    assign inter_8[546] = inter_7[546]^inter_7[674];
    assign inter_8[547] = inter_7[547]^inter_7[675];
    assign inter_8[548] = inter_7[548]^inter_7[676];
    assign inter_8[549] = inter_7[549]^inter_7[677];
    assign inter_8[550] = inter_7[550]^inter_7[678];
    assign inter_8[551] = inter_7[551]^inter_7[679];
    assign inter_8[552] = inter_7[552]^inter_7[680];
    assign inter_8[553] = inter_7[553]^inter_7[681];
    assign inter_8[554] = inter_7[554]^inter_7[682];
    assign inter_8[555] = inter_7[555]^inter_7[683];
    assign inter_8[556] = inter_7[556]^inter_7[684];
    assign inter_8[557] = inter_7[557]^inter_7[685];
    assign inter_8[558] = inter_7[558]^inter_7[686];
    assign inter_8[559] = inter_7[559]^inter_7[687];
    assign inter_8[560] = inter_7[560]^inter_7[688];
    assign inter_8[561] = inter_7[561]^inter_7[689];
    assign inter_8[562] = inter_7[562]^inter_7[690];
    assign inter_8[563] = inter_7[563]^inter_7[691];
    assign inter_8[564] = inter_7[564]^inter_7[692];
    assign inter_8[565] = inter_7[565]^inter_7[693];
    assign inter_8[566] = inter_7[566]^inter_7[694];
    assign inter_8[567] = inter_7[567]^inter_7[695];
    assign inter_8[568] = inter_7[568]^inter_7[696];
    assign inter_8[569] = inter_7[569]^inter_7[697];
    assign inter_8[570] = inter_7[570]^inter_7[698];
    assign inter_8[571] = inter_7[571]^inter_7[699];
    assign inter_8[572] = inter_7[572]^inter_7[700];
    assign inter_8[573] = inter_7[573]^inter_7[701];
    assign inter_8[574] = inter_7[574]^inter_7[702];
    assign inter_8[575] = inter_7[575]^inter_7[703];
    assign inter_8[576] = inter_7[576]^inter_7[704];
    assign inter_8[577] = inter_7[577]^inter_7[705];
    assign inter_8[578] = inter_7[578]^inter_7[706];
    assign inter_8[579] = inter_7[579]^inter_7[707];
    assign inter_8[580] = inter_7[580]^inter_7[708];
    assign inter_8[581] = inter_7[581]^inter_7[709];
    assign inter_8[582] = inter_7[582]^inter_7[710];
    assign inter_8[583] = inter_7[583]^inter_7[711];
    assign inter_8[584] = inter_7[584]^inter_7[712];
    assign inter_8[585] = inter_7[585]^inter_7[713];
    assign inter_8[586] = inter_7[586]^inter_7[714];
    assign inter_8[587] = inter_7[587]^inter_7[715];
    assign inter_8[588] = inter_7[588]^inter_7[716];
    assign inter_8[589] = inter_7[589]^inter_7[717];
    assign inter_8[590] = inter_7[590]^inter_7[718];
    assign inter_8[591] = inter_7[591]^inter_7[719];
    assign inter_8[592] = inter_7[592]^inter_7[720];
    assign inter_8[593] = inter_7[593]^inter_7[721];
    assign inter_8[594] = inter_7[594]^inter_7[722];
    assign inter_8[595] = inter_7[595]^inter_7[723];
    assign inter_8[596] = inter_7[596]^inter_7[724];
    assign inter_8[597] = inter_7[597]^inter_7[725];
    assign inter_8[598] = inter_7[598]^inter_7[726];
    assign inter_8[599] = inter_7[599]^inter_7[727];
    assign inter_8[600] = inter_7[600]^inter_7[728];
    assign inter_8[601] = inter_7[601]^inter_7[729];
    assign inter_8[602] = inter_7[602]^inter_7[730];
    assign inter_8[603] = inter_7[603]^inter_7[731];
    assign inter_8[604] = inter_7[604]^inter_7[732];
    assign inter_8[605] = inter_7[605]^inter_7[733];
    assign inter_8[606] = inter_7[606]^inter_7[734];
    assign inter_8[607] = inter_7[607]^inter_7[735];
    assign inter_8[608] = inter_7[608]^inter_7[736];
    assign inter_8[609] = inter_7[609]^inter_7[737];
    assign inter_8[610] = inter_7[610]^inter_7[738];
    assign inter_8[611] = inter_7[611]^inter_7[739];
    assign inter_8[612] = inter_7[612]^inter_7[740];
    assign inter_8[613] = inter_7[613]^inter_7[741];
    assign inter_8[614] = inter_7[614]^inter_7[742];
    assign inter_8[615] = inter_7[615]^inter_7[743];
    assign inter_8[616] = inter_7[616]^inter_7[744];
    assign inter_8[617] = inter_7[617]^inter_7[745];
    assign inter_8[618] = inter_7[618]^inter_7[746];
    assign inter_8[619] = inter_7[619]^inter_7[747];
    assign inter_8[620] = inter_7[620]^inter_7[748];
    assign inter_8[621] = inter_7[621]^inter_7[749];
    assign inter_8[622] = inter_7[622]^inter_7[750];
    assign inter_8[623] = inter_7[623]^inter_7[751];
    assign inter_8[624] = inter_7[624]^inter_7[752];
    assign inter_8[625] = inter_7[625]^inter_7[753];
    assign inter_8[626] = inter_7[626]^inter_7[754];
    assign inter_8[627] = inter_7[627]^inter_7[755];
    assign inter_8[628] = inter_7[628]^inter_7[756];
    assign inter_8[629] = inter_7[629]^inter_7[757];
    assign inter_8[630] = inter_7[630]^inter_7[758];
    assign inter_8[631] = inter_7[631]^inter_7[759];
    assign inter_8[632] = inter_7[632]^inter_7[760];
    assign inter_8[633] = inter_7[633]^inter_7[761];
    assign inter_8[634] = inter_7[634]^inter_7[762];
    assign inter_8[635] = inter_7[635]^inter_7[763];
    assign inter_8[636] = inter_7[636]^inter_7[764];
    assign inter_8[637] = inter_7[637]^inter_7[765];
    assign inter_8[638] = inter_7[638]^inter_7[766];
    assign inter_8[639] = inter_7[639]^inter_7[767];
    assign inter_8[640] = inter_7[640];
    assign inter_8[641] = inter_7[641];
    assign inter_8[642] = inter_7[642];
    assign inter_8[643] = inter_7[643];
    assign inter_8[644] = inter_7[644];
    assign inter_8[645] = inter_7[645];
    assign inter_8[646] = inter_7[646];
    assign inter_8[647] = inter_7[647];
    assign inter_8[648] = inter_7[648];
    assign inter_8[649] = inter_7[649];
    assign inter_8[650] = inter_7[650];
    assign inter_8[651] = inter_7[651];
    assign inter_8[652] = inter_7[652];
    assign inter_8[653] = inter_7[653];
    assign inter_8[654] = inter_7[654];
    assign inter_8[655] = inter_7[655];
    assign inter_8[656] = inter_7[656];
    assign inter_8[657] = inter_7[657];
    assign inter_8[658] = inter_7[658];
    assign inter_8[659] = inter_7[659];
    assign inter_8[660] = inter_7[660];
    assign inter_8[661] = inter_7[661];
    assign inter_8[662] = inter_7[662];
    assign inter_8[663] = inter_7[663];
    assign inter_8[664] = inter_7[664];
    assign inter_8[665] = inter_7[665];
    assign inter_8[666] = inter_7[666];
    assign inter_8[667] = inter_7[667];
    assign inter_8[668] = inter_7[668];
    assign inter_8[669] = inter_7[669];
    assign inter_8[670] = inter_7[670];
    assign inter_8[671] = inter_7[671];
    assign inter_8[672] = inter_7[672];
    assign inter_8[673] = inter_7[673];
    assign inter_8[674] = inter_7[674];
    assign inter_8[675] = inter_7[675];
    assign inter_8[676] = inter_7[676];
    assign inter_8[677] = inter_7[677];
    assign inter_8[678] = inter_7[678];
    assign inter_8[679] = inter_7[679];
    assign inter_8[680] = inter_7[680];
    assign inter_8[681] = inter_7[681];
    assign inter_8[682] = inter_7[682];
    assign inter_8[683] = inter_7[683];
    assign inter_8[684] = inter_7[684];
    assign inter_8[685] = inter_7[685];
    assign inter_8[686] = inter_7[686];
    assign inter_8[687] = inter_7[687];
    assign inter_8[688] = inter_7[688];
    assign inter_8[689] = inter_7[689];
    assign inter_8[690] = inter_7[690];
    assign inter_8[691] = inter_7[691];
    assign inter_8[692] = inter_7[692];
    assign inter_8[693] = inter_7[693];
    assign inter_8[694] = inter_7[694];
    assign inter_8[695] = inter_7[695];
    assign inter_8[696] = inter_7[696];
    assign inter_8[697] = inter_7[697];
    assign inter_8[698] = inter_7[698];
    assign inter_8[699] = inter_7[699];
    assign inter_8[700] = inter_7[700];
    assign inter_8[701] = inter_7[701];
    assign inter_8[702] = inter_7[702];
    assign inter_8[703] = inter_7[703];
    assign inter_8[704] = inter_7[704];
    assign inter_8[705] = inter_7[705];
    assign inter_8[706] = inter_7[706];
    assign inter_8[707] = inter_7[707];
    assign inter_8[708] = inter_7[708];
    assign inter_8[709] = inter_7[709];
    assign inter_8[710] = inter_7[710];
    assign inter_8[711] = inter_7[711];
    assign inter_8[712] = inter_7[712];
    assign inter_8[713] = inter_7[713];
    assign inter_8[714] = inter_7[714];
    assign inter_8[715] = inter_7[715];
    assign inter_8[716] = inter_7[716];
    assign inter_8[717] = inter_7[717];
    assign inter_8[718] = inter_7[718];
    assign inter_8[719] = inter_7[719];
    assign inter_8[720] = inter_7[720];
    assign inter_8[721] = inter_7[721];
    assign inter_8[722] = inter_7[722];
    assign inter_8[723] = inter_7[723];
    assign inter_8[724] = inter_7[724];
    assign inter_8[725] = inter_7[725];
    assign inter_8[726] = inter_7[726];
    assign inter_8[727] = inter_7[727];
    assign inter_8[728] = inter_7[728];
    assign inter_8[729] = inter_7[729];
    assign inter_8[730] = inter_7[730];
    assign inter_8[731] = inter_7[731];
    assign inter_8[732] = inter_7[732];
    assign inter_8[733] = inter_7[733];
    assign inter_8[734] = inter_7[734];
    assign inter_8[735] = inter_7[735];
    assign inter_8[736] = inter_7[736];
    assign inter_8[737] = inter_7[737];
    assign inter_8[738] = inter_7[738];
    assign inter_8[739] = inter_7[739];
    assign inter_8[740] = inter_7[740];
    assign inter_8[741] = inter_7[741];
    assign inter_8[742] = inter_7[742];
    assign inter_8[743] = inter_7[743];
    assign inter_8[744] = inter_7[744];
    assign inter_8[745] = inter_7[745];
    assign inter_8[746] = inter_7[746];
    assign inter_8[747] = inter_7[747];
    assign inter_8[748] = inter_7[748];
    assign inter_8[749] = inter_7[749];
    assign inter_8[750] = inter_7[750];
    assign inter_8[751] = inter_7[751];
    assign inter_8[752] = inter_7[752];
    assign inter_8[753] = inter_7[753];
    assign inter_8[754] = inter_7[754];
    assign inter_8[755] = inter_7[755];
    assign inter_8[756] = inter_7[756];
    assign inter_8[757] = inter_7[757];
    assign inter_8[758] = inter_7[758];
    assign inter_8[759] = inter_7[759];
    assign inter_8[760] = inter_7[760];
    assign inter_8[761] = inter_7[761];
    assign inter_8[762] = inter_7[762];
    assign inter_8[763] = inter_7[763];
    assign inter_8[764] = inter_7[764];
    assign inter_8[765] = inter_7[765];
    assign inter_8[766] = inter_7[766];
    assign inter_8[767] = inter_7[767];
    assign inter_8[768] = inter_7[768]^inter_7[896];
    assign inter_8[769] = inter_7[769]^inter_7[897];
    assign inter_8[770] = inter_7[770]^inter_7[898];
    assign inter_8[771] = inter_7[771]^inter_7[899];
    assign inter_8[772] = inter_7[772]^inter_7[900];
    assign inter_8[773] = inter_7[773]^inter_7[901];
    assign inter_8[774] = inter_7[774]^inter_7[902];
    assign inter_8[775] = inter_7[775]^inter_7[903];
    assign inter_8[776] = inter_7[776]^inter_7[904];
    assign inter_8[777] = inter_7[777]^inter_7[905];
    assign inter_8[778] = inter_7[778]^inter_7[906];
    assign inter_8[779] = inter_7[779]^inter_7[907];
    assign inter_8[780] = inter_7[780]^inter_7[908];
    assign inter_8[781] = inter_7[781]^inter_7[909];
    assign inter_8[782] = inter_7[782]^inter_7[910];
    assign inter_8[783] = inter_7[783]^inter_7[911];
    assign inter_8[784] = inter_7[784]^inter_7[912];
    assign inter_8[785] = inter_7[785]^inter_7[913];
    assign inter_8[786] = inter_7[786]^inter_7[914];
    assign inter_8[787] = inter_7[787]^inter_7[915];
    assign inter_8[788] = inter_7[788]^inter_7[916];
    assign inter_8[789] = inter_7[789]^inter_7[917];
    assign inter_8[790] = inter_7[790]^inter_7[918];
    assign inter_8[791] = inter_7[791]^inter_7[919];
    assign inter_8[792] = inter_7[792]^inter_7[920];
    assign inter_8[793] = inter_7[793]^inter_7[921];
    assign inter_8[794] = inter_7[794]^inter_7[922];
    assign inter_8[795] = inter_7[795]^inter_7[923];
    assign inter_8[796] = inter_7[796]^inter_7[924];
    assign inter_8[797] = inter_7[797]^inter_7[925];
    assign inter_8[798] = inter_7[798]^inter_7[926];
    assign inter_8[799] = inter_7[799]^inter_7[927];
    assign inter_8[800] = inter_7[800]^inter_7[928];
    assign inter_8[801] = inter_7[801]^inter_7[929];
    assign inter_8[802] = inter_7[802]^inter_7[930];
    assign inter_8[803] = inter_7[803]^inter_7[931];
    assign inter_8[804] = inter_7[804]^inter_7[932];
    assign inter_8[805] = inter_7[805]^inter_7[933];
    assign inter_8[806] = inter_7[806]^inter_7[934];
    assign inter_8[807] = inter_7[807]^inter_7[935];
    assign inter_8[808] = inter_7[808]^inter_7[936];
    assign inter_8[809] = inter_7[809]^inter_7[937];
    assign inter_8[810] = inter_7[810]^inter_7[938];
    assign inter_8[811] = inter_7[811]^inter_7[939];
    assign inter_8[812] = inter_7[812]^inter_7[940];
    assign inter_8[813] = inter_7[813]^inter_7[941];
    assign inter_8[814] = inter_7[814]^inter_7[942];
    assign inter_8[815] = inter_7[815]^inter_7[943];
    assign inter_8[816] = inter_7[816]^inter_7[944];
    assign inter_8[817] = inter_7[817]^inter_7[945];
    assign inter_8[818] = inter_7[818]^inter_7[946];
    assign inter_8[819] = inter_7[819]^inter_7[947];
    assign inter_8[820] = inter_7[820]^inter_7[948];
    assign inter_8[821] = inter_7[821]^inter_7[949];
    assign inter_8[822] = inter_7[822]^inter_7[950];
    assign inter_8[823] = inter_7[823]^inter_7[951];
    assign inter_8[824] = inter_7[824]^inter_7[952];
    assign inter_8[825] = inter_7[825]^inter_7[953];
    assign inter_8[826] = inter_7[826]^inter_7[954];
    assign inter_8[827] = inter_7[827]^inter_7[955];
    assign inter_8[828] = inter_7[828]^inter_7[956];
    assign inter_8[829] = inter_7[829]^inter_7[957];
    assign inter_8[830] = inter_7[830]^inter_7[958];
    assign inter_8[831] = inter_7[831]^inter_7[959];
    assign inter_8[832] = inter_7[832]^inter_7[960];
    assign inter_8[833] = inter_7[833]^inter_7[961];
    assign inter_8[834] = inter_7[834]^inter_7[962];
    assign inter_8[835] = inter_7[835]^inter_7[963];
    assign inter_8[836] = inter_7[836]^inter_7[964];
    assign inter_8[837] = inter_7[837]^inter_7[965];
    assign inter_8[838] = inter_7[838]^inter_7[966];
    assign inter_8[839] = inter_7[839]^inter_7[967];
    assign inter_8[840] = inter_7[840]^inter_7[968];
    assign inter_8[841] = inter_7[841]^inter_7[969];
    assign inter_8[842] = inter_7[842]^inter_7[970];
    assign inter_8[843] = inter_7[843]^inter_7[971];
    assign inter_8[844] = inter_7[844]^inter_7[972];
    assign inter_8[845] = inter_7[845]^inter_7[973];
    assign inter_8[846] = inter_7[846]^inter_7[974];
    assign inter_8[847] = inter_7[847]^inter_7[975];
    assign inter_8[848] = inter_7[848]^inter_7[976];
    assign inter_8[849] = inter_7[849]^inter_7[977];
    assign inter_8[850] = inter_7[850]^inter_7[978];
    assign inter_8[851] = inter_7[851]^inter_7[979];
    assign inter_8[852] = inter_7[852]^inter_7[980];
    assign inter_8[853] = inter_7[853]^inter_7[981];
    assign inter_8[854] = inter_7[854]^inter_7[982];
    assign inter_8[855] = inter_7[855]^inter_7[983];
    assign inter_8[856] = inter_7[856]^inter_7[984];
    assign inter_8[857] = inter_7[857]^inter_7[985];
    assign inter_8[858] = inter_7[858]^inter_7[986];
    assign inter_8[859] = inter_7[859]^inter_7[987];
    assign inter_8[860] = inter_7[860]^inter_7[988];
    assign inter_8[861] = inter_7[861]^inter_7[989];
    assign inter_8[862] = inter_7[862]^inter_7[990];
    assign inter_8[863] = inter_7[863]^inter_7[991];
    assign inter_8[864] = inter_7[864]^inter_7[992];
    assign inter_8[865] = inter_7[865]^inter_7[993];
    assign inter_8[866] = inter_7[866]^inter_7[994];
    assign inter_8[867] = inter_7[867]^inter_7[995];
    assign inter_8[868] = inter_7[868]^inter_7[996];
    assign inter_8[869] = inter_7[869]^inter_7[997];
    assign inter_8[870] = inter_7[870]^inter_7[998];
    assign inter_8[871] = inter_7[871]^inter_7[999];
    assign inter_8[872] = inter_7[872]^inter_7[1000];
    assign inter_8[873] = inter_7[873]^inter_7[1001];
    assign inter_8[874] = inter_7[874]^inter_7[1002];
    assign inter_8[875] = inter_7[875]^inter_7[1003];
    assign inter_8[876] = inter_7[876]^inter_7[1004];
    assign inter_8[877] = inter_7[877]^inter_7[1005];
    assign inter_8[878] = inter_7[878]^inter_7[1006];
    assign inter_8[879] = inter_7[879]^inter_7[1007];
    assign inter_8[880] = inter_7[880]^inter_7[1008];
    assign inter_8[881] = inter_7[881]^inter_7[1009];
    assign inter_8[882] = inter_7[882]^inter_7[1010];
    assign inter_8[883] = inter_7[883]^inter_7[1011];
    assign inter_8[884] = inter_7[884]^inter_7[1012];
    assign inter_8[885] = inter_7[885]^inter_7[1013];
    assign inter_8[886] = inter_7[886]^inter_7[1014];
    assign inter_8[887] = inter_7[887]^inter_7[1015];
    assign inter_8[888] = inter_7[888]^inter_7[1016];
    assign inter_8[889] = inter_7[889]^inter_7[1017];
    assign inter_8[890] = inter_7[890]^inter_7[1018];
    assign inter_8[891] = inter_7[891]^inter_7[1019];
    assign inter_8[892] = inter_7[892]^inter_7[1020];
    assign inter_8[893] = inter_7[893]^inter_7[1021];
    assign inter_8[894] = inter_7[894]^inter_7[1022];
    assign inter_8[895] = inter_7[895]^inter_7[1023];
    assign inter_8[896] = inter_7[896];
    assign inter_8[897] = inter_7[897];
    assign inter_8[898] = inter_7[898];
    assign inter_8[899] = inter_7[899];
    assign inter_8[900] = inter_7[900];
    assign inter_8[901] = inter_7[901];
    assign inter_8[902] = inter_7[902];
    assign inter_8[903] = inter_7[903];
    assign inter_8[904] = inter_7[904];
    assign inter_8[905] = inter_7[905];
    assign inter_8[906] = inter_7[906];
    assign inter_8[907] = inter_7[907];
    assign inter_8[908] = inter_7[908];
    assign inter_8[909] = inter_7[909];
    assign inter_8[910] = inter_7[910];
    assign inter_8[911] = inter_7[911];
    assign inter_8[912] = inter_7[912];
    assign inter_8[913] = inter_7[913];
    assign inter_8[914] = inter_7[914];
    assign inter_8[915] = inter_7[915];
    assign inter_8[916] = inter_7[916];
    assign inter_8[917] = inter_7[917];
    assign inter_8[918] = inter_7[918];
    assign inter_8[919] = inter_7[919];
    assign inter_8[920] = inter_7[920];
    assign inter_8[921] = inter_7[921];
    assign inter_8[922] = inter_7[922];
    assign inter_8[923] = inter_7[923];
    assign inter_8[924] = inter_7[924];
    assign inter_8[925] = inter_7[925];
    assign inter_8[926] = inter_7[926];
    assign inter_8[927] = inter_7[927];
    assign inter_8[928] = inter_7[928];
    assign inter_8[929] = inter_7[929];
    assign inter_8[930] = inter_7[930];
    assign inter_8[931] = inter_7[931];
    assign inter_8[932] = inter_7[932];
    assign inter_8[933] = inter_7[933];
    assign inter_8[934] = inter_7[934];
    assign inter_8[935] = inter_7[935];
    assign inter_8[936] = inter_7[936];
    assign inter_8[937] = inter_7[937];
    assign inter_8[938] = inter_7[938];
    assign inter_8[939] = inter_7[939];
    assign inter_8[940] = inter_7[940];
    assign inter_8[941] = inter_7[941];
    assign inter_8[942] = inter_7[942];
    assign inter_8[943] = inter_7[943];
    assign inter_8[944] = inter_7[944];
    assign inter_8[945] = inter_7[945];
    assign inter_8[946] = inter_7[946];
    assign inter_8[947] = inter_7[947];
    assign inter_8[948] = inter_7[948];
    assign inter_8[949] = inter_7[949];
    assign inter_8[950] = inter_7[950];
    assign inter_8[951] = inter_7[951];
    assign inter_8[952] = inter_7[952];
    assign inter_8[953] = inter_7[953];
    assign inter_8[954] = inter_7[954];
    assign inter_8[955] = inter_7[955];
    assign inter_8[956] = inter_7[956];
    assign inter_8[957] = inter_7[957];
    assign inter_8[958] = inter_7[958];
    assign inter_8[959] = inter_7[959];
    assign inter_8[960] = inter_7[960];
    assign inter_8[961] = inter_7[961];
    assign inter_8[962] = inter_7[962];
    assign inter_8[963] = inter_7[963];
    assign inter_8[964] = inter_7[964];
    assign inter_8[965] = inter_7[965];
    assign inter_8[966] = inter_7[966];
    assign inter_8[967] = inter_7[967];
    assign inter_8[968] = inter_7[968];
    assign inter_8[969] = inter_7[969];
    assign inter_8[970] = inter_7[970];
    assign inter_8[971] = inter_7[971];
    assign inter_8[972] = inter_7[972];
    assign inter_8[973] = inter_7[973];
    assign inter_8[974] = inter_7[974];
    assign inter_8[975] = inter_7[975];
    assign inter_8[976] = inter_7[976];
    assign inter_8[977] = inter_7[977];
    assign inter_8[978] = inter_7[978];
    assign inter_8[979] = inter_7[979];
    assign inter_8[980] = inter_7[980];
    assign inter_8[981] = inter_7[981];
    assign inter_8[982] = inter_7[982];
    assign inter_8[983] = inter_7[983];
    assign inter_8[984] = inter_7[984];
    assign inter_8[985] = inter_7[985];
    assign inter_8[986] = inter_7[986];
    assign inter_8[987] = inter_7[987];
    assign inter_8[988] = inter_7[988];
    assign inter_8[989] = inter_7[989];
    assign inter_8[990] = inter_7[990];
    assign inter_8[991] = inter_7[991];
    assign inter_8[992] = inter_7[992];
    assign inter_8[993] = inter_7[993];
    assign inter_8[994] = inter_7[994];
    assign inter_8[995] = inter_7[995];
    assign inter_8[996] = inter_7[996];
    assign inter_8[997] = inter_7[997];
    assign inter_8[998] = inter_7[998];
    assign inter_8[999] = inter_7[999];
    assign inter_8[1000] = inter_7[1000];
    assign inter_8[1001] = inter_7[1001];
    assign inter_8[1002] = inter_7[1002];
    assign inter_8[1003] = inter_7[1003];
    assign inter_8[1004] = inter_7[1004];
    assign inter_8[1005] = inter_7[1005];
    assign inter_8[1006] = inter_7[1006];
    assign inter_8[1007] = inter_7[1007];
    assign inter_8[1008] = inter_7[1008];
    assign inter_8[1009] = inter_7[1009];
    assign inter_8[1010] = inter_7[1010];
    assign inter_8[1011] = inter_7[1011];
    assign inter_8[1012] = inter_7[1012];
    assign inter_8[1013] = inter_7[1013];
    assign inter_8[1014] = inter_7[1014];
    assign inter_8[1015] = inter_7[1015];
    assign inter_8[1016] = inter_7[1016];
    assign inter_8[1017] = inter_7[1017];
    assign inter_8[1018] = inter_7[1018];
    assign inter_8[1019] = inter_7[1019];
    assign inter_8[1020] = inter_7[1020];
    assign inter_8[1021] = inter_7[1021];
    assign inter_8[1022] = inter_7[1022];
    assign inter_8[1023] = inter_7[1023];
    /***************************/
    assign inter_9[0] = inter_8[0]^inter_8[256];
    assign inter_9[1] = inter_8[1]^inter_8[257];
    assign inter_9[2] = inter_8[2]^inter_8[258];
    assign inter_9[3] = inter_8[3]^inter_8[259];
    assign inter_9[4] = inter_8[4]^inter_8[260];
    assign inter_9[5] = inter_8[5]^inter_8[261];
    assign inter_9[6] = inter_8[6]^inter_8[262];
    assign inter_9[7] = inter_8[7]^inter_8[263];
    assign inter_9[8] = inter_8[8]^inter_8[264];
    assign inter_9[9] = inter_8[9]^inter_8[265];
    assign inter_9[10] = inter_8[10]^inter_8[266];
    assign inter_9[11] = inter_8[11]^inter_8[267];
    assign inter_9[12] = inter_8[12]^inter_8[268];
    assign inter_9[13] = inter_8[13]^inter_8[269];
    assign inter_9[14] = inter_8[14]^inter_8[270];
    assign inter_9[15] = inter_8[15]^inter_8[271];
    assign inter_9[16] = inter_8[16]^inter_8[272];
    assign inter_9[17] = inter_8[17]^inter_8[273];
    assign inter_9[18] = inter_8[18]^inter_8[274];
    assign inter_9[19] = inter_8[19]^inter_8[275];
    assign inter_9[20] = inter_8[20]^inter_8[276];
    assign inter_9[21] = inter_8[21]^inter_8[277];
    assign inter_9[22] = inter_8[22]^inter_8[278];
    assign inter_9[23] = inter_8[23]^inter_8[279];
    assign inter_9[24] = inter_8[24]^inter_8[280];
    assign inter_9[25] = inter_8[25]^inter_8[281];
    assign inter_9[26] = inter_8[26]^inter_8[282];
    assign inter_9[27] = inter_8[27]^inter_8[283];
    assign inter_9[28] = inter_8[28]^inter_8[284];
    assign inter_9[29] = inter_8[29]^inter_8[285];
    assign inter_9[30] = inter_8[30]^inter_8[286];
    assign inter_9[31] = inter_8[31]^inter_8[287];
    assign inter_9[32] = inter_8[32]^inter_8[288];
    assign inter_9[33] = inter_8[33]^inter_8[289];
    assign inter_9[34] = inter_8[34]^inter_8[290];
    assign inter_9[35] = inter_8[35]^inter_8[291];
    assign inter_9[36] = inter_8[36]^inter_8[292];
    assign inter_9[37] = inter_8[37]^inter_8[293];
    assign inter_9[38] = inter_8[38]^inter_8[294];
    assign inter_9[39] = inter_8[39]^inter_8[295];
    assign inter_9[40] = inter_8[40]^inter_8[296];
    assign inter_9[41] = inter_8[41]^inter_8[297];
    assign inter_9[42] = inter_8[42]^inter_8[298];
    assign inter_9[43] = inter_8[43]^inter_8[299];
    assign inter_9[44] = inter_8[44]^inter_8[300];
    assign inter_9[45] = inter_8[45]^inter_8[301];
    assign inter_9[46] = inter_8[46]^inter_8[302];
    assign inter_9[47] = inter_8[47]^inter_8[303];
    assign inter_9[48] = inter_8[48]^inter_8[304];
    assign inter_9[49] = inter_8[49]^inter_8[305];
    assign inter_9[50] = inter_8[50]^inter_8[306];
    assign inter_9[51] = inter_8[51]^inter_8[307];
    assign inter_9[52] = inter_8[52]^inter_8[308];
    assign inter_9[53] = inter_8[53]^inter_8[309];
    assign inter_9[54] = inter_8[54]^inter_8[310];
    assign inter_9[55] = inter_8[55]^inter_8[311];
    assign inter_9[56] = inter_8[56]^inter_8[312];
    assign inter_9[57] = inter_8[57]^inter_8[313];
    assign inter_9[58] = inter_8[58]^inter_8[314];
    assign inter_9[59] = inter_8[59]^inter_8[315];
    assign inter_9[60] = inter_8[60]^inter_8[316];
    assign inter_9[61] = inter_8[61]^inter_8[317];
    assign inter_9[62] = inter_8[62]^inter_8[318];
    assign inter_9[63] = inter_8[63]^inter_8[319];
    assign inter_9[64] = inter_8[64]^inter_8[320];
    assign inter_9[65] = inter_8[65]^inter_8[321];
    assign inter_9[66] = inter_8[66]^inter_8[322];
    assign inter_9[67] = inter_8[67]^inter_8[323];
    assign inter_9[68] = inter_8[68]^inter_8[324];
    assign inter_9[69] = inter_8[69]^inter_8[325];
    assign inter_9[70] = inter_8[70]^inter_8[326];
    assign inter_9[71] = inter_8[71]^inter_8[327];
    assign inter_9[72] = inter_8[72]^inter_8[328];
    assign inter_9[73] = inter_8[73]^inter_8[329];
    assign inter_9[74] = inter_8[74]^inter_8[330];
    assign inter_9[75] = inter_8[75]^inter_8[331];
    assign inter_9[76] = inter_8[76]^inter_8[332];
    assign inter_9[77] = inter_8[77]^inter_8[333];
    assign inter_9[78] = inter_8[78]^inter_8[334];
    assign inter_9[79] = inter_8[79]^inter_8[335];
    assign inter_9[80] = inter_8[80]^inter_8[336];
    assign inter_9[81] = inter_8[81]^inter_8[337];
    assign inter_9[82] = inter_8[82]^inter_8[338];
    assign inter_9[83] = inter_8[83]^inter_8[339];
    assign inter_9[84] = inter_8[84]^inter_8[340];
    assign inter_9[85] = inter_8[85]^inter_8[341];
    assign inter_9[86] = inter_8[86]^inter_8[342];
    assign inter_9[87] = inter_8[87]^inter_8[343];
    assign inter_9[88] = inter_8[88]^inter_8[344];
    assign inter_9[89] = inter_8[89]^inter_8[345];
    assign inter_9[90] = inter_8[90]^inter_8[346];
    assign inter_9[91] = inter_8[91]^inter_8[347];
    assign inter_9[92] = inter_8[92]^inter_8[348];
    assign inter_9[93] = inter_8[93]^inter_8[349];
    assign inter_9[94] = inter_8[94]^inter_8[350];
    assign inter_9[95] = inter_8[95]^inter_8[351];
    assign inter_9[96] = inter_8[96]^inter_8[352];
    assign inter_9[97] = inter_8[97]^inter_8[353];
    assign inter_9[98] = inter_8[98]^inter_8[354];
    assign inter_9[99] = inter_8[99]^inter_8[355];
    assign inter_9[100] = inter_8[100]^inter_8[356];
    assign inter_9[101] = inter_8[101]^inter_8[357];
    assign inter_9[102] = inter_8[102]^inter_8[358];
    assign inter_9[103] = inter_8[103]^inter_8[359];
    assign inter_9[104] = inter_8[104]^inter_8[360];
    assign inter_9[105] = inter_8[105]^inter_8[361];
    assign inter_9[106] = inter_8[106]^inter_8[362];
    assign inter_9[107] = inter_8[107]^inter_8[363];
    assign inter_9[108] = inter_8[108]^inter_8[364];
    assign inter_9[109] = inter_8[109]^inter_8[365];
    assign inter_9[110] = inter_8[110]^inter_8[366];
    assign inter_9[111] = inter_8[111]^inter_8[367];
    assign inter_9[112] = inter_8[112]^inter_8[368];
    assign inter_9[113] = inter_8[113]^inter_8[369];
    assign inter_9[114] = inter_8[114]^inter_8[370];
    assign inter_9[115] = inter_8[115]^inter_8[371];
    assign inter_9[116] = inter_8[116]^inter_8[372];
    assign inter_9[117] = inter_8[117]^inter_8[373];
    assign inter_9[118] = inter_8[118]^inter_8[374];
    assign inter_9[119] = inter_8[119]^inter_8[375];
    assign inter_9[120] = inter_8[120]^inter_8[376];
    assign inter_9[121] = inter_8[121]^inter_8[377];
    assign inter_9[122] = inter_8[122]^inter_8[378];
    assign inter_9[123] = inter_8[123]^inter_8[379];
    assign inter_9[124] = inter_8[124]^inter_8[380];
    assign inter_9[125] = inter_8[125]^inter_8[381];
    assign inter_9[126] = inter_8[126]^inter_8[382];
    assign inter_9[127] = inter_8[127]^inter_8[383];
    assign inter_9[128] = inter_8[128]^inter_8[384];
    assign inter_9[129] = inter_8[129]^inter_8[385];
    assign inter_9[130] = inter_8[130]^inter_8[386];
    assign inter_9[131] = inter_8[131]^inter_8[387];
    assign inter_9[132] = inter_8[132]^inter_8[388];
    assign inter_9[133] = inter_8[133]^inter_8[389];
    assign inter_9[134] = inter_8[134]^inter_8[390];
    assign inter_9[135] = inter_8[135]^inter_8[391];
    assign inter_9[136] = inter_8[136]^inter_8[392];
    assign inter_9[137] = inter_8[137]^inter_8[393];
    assign inter_9[138] = inter_8[138]^inter_8[394];
    assign inter_9[139] = inter_8[139]^inter_8[395];
    assign inter_9[140] = inter_8[140]^inter_8[396];
    assign inter_9[141] = inter_8[141]^inter_8[397];
    assign inter_9[142] = inter_8[142]^inter_8[398];
    assign inter_9[143] = inter_8[143]^inter_8[399];
    assign inter_9[144] = inter_8[144]^inter_8[400];
    assign inter_9[145] = inter_8[145]^inter_8[401];
    assign inter_9[146] = inter_8[146]^inter_8[402];
    assign inter_9[147] = inter_8[147]^inter_8[403];
    assign inter_9[148] = inter_8[148]^inter_8[404];
    assign inter_9[149] = inter_8[149]^inter_8[405];
    assign inter_9[150] = inter_8[150]^inter_8[406];
    assign inter_9[151] = inter_8[151]^inter_8[407];
    assign inter_9[152] = inter_8[152]^inter_8[408];
    assign inter_9[153] = inter_8[153]^inter_8[409];
    assign inter_9[154] = inter_8[154]^inter_8[410];
    assign inter_9[155] = inter_8[155]^inter_8[411];
    assign inter_9[156] = inter_8[156]^inter_8[412];
    assign inter_9[157] = inter_8[157]^inter_8[413];
    assign inter_9[158] = inter_8[158]^inter_8[414];
    assign inter_9[159] = inter_8[159]^inter_8[415];
    assign inter_9[160] = inter_8[160]^inter_8[416];
    assign inter_9[161] = inter_8[161]^inter_8[417];
    assign inter_9[162] = inter_8[162]^inter_8[418];
    assign inter_9[163] = inter_8[163]^inter_8[419];
    assign inter_9[164] = inter_8[164]^inter_8[420];
    assign inter_9[165] = inter_8[165]^inter_8[421];
    assign inter_9[166] = inter_8[166]^inter_8[422];
    assign inter_9[167] = inter_8[167]^inter_8[423];
    assign inter_9[168] = inter_8[168]^inter_8[424];
    assign inter_9[169] = inter_8[169]^inter_8[425];
    assign inter_9[170] = inter_8[170]^inter_8[426];
    assign inter_9[171] = inter_8[171]^inter_8[427];
    assign inter_9[172] = inter_8[172]^inter_8[428];
    assign inter_9[173] = inter_8[173]^inter_8[429];
    assign inter_9[174] = inter_8[174]^inter_8[430];
    assign inter_9[175] = inter_8[175]^inter_8[431];
    assign inter_9[176] = inter_8[176]^inter_8[432];
    assign inter_9[177] = inter_8[177]^inter_8[433];
    assign inter_9[178] = inter_8[178]^inter_8[434];
    assign inter_9[179] = inter_8[179]^inter_8[435];
    assign inter_9[180] = inter_8[180]^inter_8[436];
    assign inter_9[181] = inter_8[181]^inter_8[437];
    assign inter_9[182] = inter_8[182]^inter_8[438];
    assign inter_9[183] = inter_8[183]^inter_8[439];
    assign inter_9[184] = inter_8[184]^inter_8[440];
    assign inter_9[185] = inter_8[185]^inter_8[441];
    assign inter_9[186] = inter_8[186]^inter_8[442];
    assign inter_9[187] = inter_8[187]^inter_8[443];
    assign inter_9[188] = inter_8[188]^inter_8[444];
    assign inter_9[189] = inter_8[189]^inter_8[445];
    assign inter_9[190] = inter_8[190]^inter_8[446];
    assign inter_9[191] = inter_8[191]^inter_8[447];
    assign inter_9[192] = inter_8[192]^inter_8[448];
    assign inter_9[193] = inter_8[193]^inter_8[449];
    assign inter_9[194] = inter_8[194]^inter_8[450];
    assign inter_9[195] = inter_8[195]^inter_8[451];
    assign inter_9[196] = inter_8[196]^inter_8[452];
    assign inter_9[197] = inter_8[197]^inter_8[453];
    assign inter_9[198] = inter_8[198]^inter_8[454];
    assign inter_9[199] = inter_8[199]^inter_8[455];
    assign inter_9[200] = inter_8[200]^inter_8[456];
    assign inter_9[201] = inter_8[201]^inter_8[457];
    assign inter_9[202] = inter_8[202]^inter_8[458];
    assign inter_9[203] = inter_8[203]^inter_8[459];
    assign inter_9[204] = inter_8[204]^inter_8[460];
    assign inter_9[205] = inter_8[205]^inter_8[461];
    assign inter_9[206] = inter_8[206]^inter_8[462];
    assign inter_9[207] = inter_8[207]^inter_8[463];
    assign inter_9[208] = inter_8[208]^inter_8[464];
    assign inter_9[209] = inter_8[209]^inter_8[465];
    assign inter_9[210] = inter_8[210]^inter_8[466];
    assign inter_9[211] = inter_8[211]^inter_8[467];
    assign inter_9[212] = inter_8[212]^inter_8[468];
    assign inter_9[213] = inter_8[213]^inter_8[469];
    assign inter_9[214] = inter_8[214]^inter_8[470];
    assign inter_9[215] = inter_8[215]^inter_8[471];
    assign inter_9[216] = inter_8[216]^inter_8[472];
    assign inter_9[217] = inter_8[217]^inter_8[473];
    assign inter_9[218] = inter_8[218]^inter_8[474];
    assign inter_9[219] = inter_8[219]^inter_8[475];
    assign inter_9[220] = inter_8[220]^inter_8[476];
    assign inter_9[221] = inter_8[221]^inter_8[477];
    assign inter_9[222] = inter_8[222]^inter_8[478];
    assign inter_9[223] = inter_8[223]^inter_8[479];
    assign inter_9[224] = inter_8[224]^inter_8[480];
    assign inter_9[225] = inter_8[225]^inter_8[481];
    assign inter_9[226] = inter_8[226]^inter_8[482];
    assign inter_9[227] = inter_8[227]^inter_8[483];
    assign inter_9[228] = inter_8[228]^inter_8[484];
    assign inter_9[229] = inter_8[229]^inter_8[485];
    assign inter_9[230] = inter_8[230]^inter_8[486];
    assign inter_9[231] = inter_8[231]^inter_8[487];
    assign inter_9[232] = inter_8[232]^inter_8[488];
    assign inter_9[233] = inter_8[233]^inter_8[489];
    assign inter_9[234] = inter_8[234]^inter_8[490];
    assign inter_9[235] = inter_8[235]^inter_8[491];
    assign inter_9[236] = inter_8[236]^inter_8[492];
    assign inter_9[237] = inter_8[237]^inter_8[493];
    assign inter_9[238] = inter_8[238]^inter_8[494];
    assign inter_9[239] = inter_8[239]^inter_8[495];
    assign inter_9[240] = inter_8[240]^inter_8[496];
    assign inter_9[241] = inter_8[241]^inter_8[497];
    assign inter_9[242] = inter_8[242]^inter_8[498];
    assign inter_9[243] = inter_8[243]^inter_8[499];
    assign inter_9[244] = inter_8[244]^inter_8[500];
    assign inter_9[245] = inter_8[245]^inter_8[501];
    assign inter_9[246] = inter_8[246]^inter_8[502];
    assign inter_9[247] = inter_8[247]^inter_8[503];
    assign inter_9[248] = inter_8[248]^inter_8[504];
    assign inter_9[249] = inter_8[249]^inter_8[505];
    assign inter_9[250] = inter_8[250]^inter_8[506];
    assign inter_9[251] = inter_8[251]^inter_8[507];
    assign inter_9[252] = inter_8[252]^inter_8[508];
    assign inter_9[253] = inter_8[253]^inter_8[509];
    assign inter_9[254] = inter_8[254]^inter_8[510];
    assign inter_9[255] = inter_8[255]^inter_8[511];
    assign inter_9[256] = inter_8[256];
    assign inter_9[257] = inter_8[257];
    assign inter_9[258] = inter_8[258];
    assign inter_9[259] = inter_8[259];
    assign inter_9[260] = inter_8[260];
    assign inter_9[261] = inter_8[261];
    assign inter_9[262] = inter_8[262];
    assign inter_9[263] = inter_8[263];
    assign inter_9[264] = inter_8[264];
    assign inter_9[265] = inter_8[265];
    assign inter_9[266] = inter_8[266];
    assign inter_9[267] = inter_8[267];
    assign inter_9[268] = inter_8[268];
    assign inter_9[269] = inter_8[269];
    assign inter_9[270] = inter_8[270];
    assign inter_9[271] = inter_8[271];
    assign inter_9[272] = inter_8[272];
    assign inter_9[273] = inter_8[273];
    assign inter_9[274] = inter_8[274];
    assign inter_9[275] = inter_8[275];
    assign inter_9[276] = inter_8[276];
    assign inter_9[277] = inter_8[277];
    assign inter_9[278] = inter_8[278];
    assign inter_9[279] = inter_8[279];
    assign inter_9[280] = inter_8[280];
    assign inter_9[281] = inter_8[281];
    assign inter_9[282] = inter_8[282];
    assign inter_9[283] = inter_8[283];
    assign inter_9[284] = inter_8[284];
    assign inter_9[285] = inter_8[285];
    assign inter_9[286] = inter_8[286];
    assign inter_9[287] = inter_8[287];
    assign inter_9[288] = inter_8[288];
    assign inter_9[289] = inter_8[289];
    assign inter_9[290] = inter_8[290];
    assign inter_9[291] = inter_8[291];
    assign inter_9[292] = inter_8[292];
    assign inter_9[293] = inter_8[293];
    assign inter_9[294] = inter_8[294];
    assign inter_9[295] = inter_8[295];
    assign inter_9[296] = inter_8[296];
    assign inter_9[297] = inter_8[297];
    assign inter_9[298] = inter_8[298];
    assign inter_9[299] = inter_8[299];
    assign inter_9[300] = inter_8[300];
    assign inter_9[301] = inter_8[301];
    assign inter_9[302] = inter_8[302];
    assign inter_9[303] = inter_8[303];
    assign inter_9[304] = inter_8[304];
    assign inter_9[305] = inter_8[305];
    assign inter_9[306] = inter_8[306];
    assign inter_9[307] = inter_8[307];
    assign inter_9[308] = inter_8[308];
    assign inter_9[309] = inter_8[309];
    assign inter_9[310] = inter_8[310];
    assign inter_9[311] = inter_8[311];
    assign inter_9[312] = inter_8[312];
    assign inter_9[313] = inter_8[313];
    assign inter_9[314] = inter_8[314];
    assign inter_9[315] = inter_8[315];
    assign inter_9[316] = inter_8[316];
    assign inter_9[317] = inter_8[317];
    assign inter_9[318] = inter_8[318];
    assign inter_9[319] = inter_8[319];
    assign inter_9[320] = inter_8[320];
    assign inter_9[321] = inter_8[321];
    assign inter_9[322] = inter_8[322];
    assign inter_9[323] = inter_8[323];
    assign inter_9[324] = inter_8[324];
    assign inter_9[325] = inter_8[325];
    assign inter_9[326] = inter_8[326];
    assign inter_9[327] = inter_8[327];
    assign inter_9[328] = inter_8[328];
    assign inter_9[329] = inter_8[329];
    assign inter_9[330] = inter_8[330];
    assign inter_9[331] = inter_8[331];
    assign inter_9[332] = inter_8[332];
    assign inter_9[333] = inter_8[333];
    assign inter_9[334] = inter_8[334];
    assign inter_9[335] = inter_8[335];
    assign inter_9[336] = inter_8[336];
    assign inter_9[337] = inter_8[337];
    assign inter_9[338] = inter_8[338];
    assign inter_9[339] = inter_8[339];
    assign inter_9[340] = inter_8[340];
    assign inter_9[341] = inter_8[341];
    assign inter_9[342] = inter_8[342];
    assign inter_9[343] = inter_8[343];
    assign inter_9[344] = inter_8[344];
    assign inter_9[345] = inter_8[345];
    assign inter_9[346] = inter_8[346];
    assign inter_9[347] = inter_8[347];
    assign inter_9[348] = inter_8[348];
    assign inter_9[349] = inter_8[349];
    assign inter_9[350] = inter_8[350];
    assign inter_9[351] = inter_8[351];
    assign inter_9[352] = inter_8[352];
    assign inter_9[353] = inter_8[353];
    assign inter_9[354] = inter_8[354];
    assign inter_9[355] = inter_8[355];
    assign inter_9[356] = inter_8[356];
    assign inter_9[357] = inter_8[357];
    assign inter_9[358] = inter_8[358];
    assign inter_9[359] = inter_8[359];
    assign inter_9[360] = inter_8[360];
    assign inter_9[361] = inter_8[361];
    assign inter_9[362] = inter_8[362];
    assign inter_9[363] = inter_8[363];
    assign inter_9[364] = inter_8[364];
    assign inter_9[365] = inter_8[365];
    assign inter_9[366] = inter_8[366];
    assign inter_9[367] = inter_8[367];
    assign inter_9[368] = inter_8[368];
    assign inter_9[369] = inter_8[369];
    assign inter_9[370] = inter_8[370];
    assign inter_9[371] = inter_8[371];
    assign inter_9[372] = inter_8[372];
    assign inter_9[373] = inter_8[373];
    assign inter_9[374] = inter_8[374];
    assign inter_9[375] = inter_8[375];
    assign inter_9[376] = inter_8[376];
    assign inter_9[377] = inter_8[377];
    assign inter_9[378] = inter_8[378];
    assign inter_9[379] = inter_8[379];
    assign inter_9[380] = inter_8[380];
    assign inter_9[381] = inter_8[381];
    assign inter_9[382] = inter_8[382];
    assign inter_9[383] = inter_8[383];
    assign inter_9[384] = inter_8[384];
    assign inter_9[385] = inter_8[385];
    assign inter_9[386] = inter_8[386];
    assign inter_9[387] = inter_8[387];
    assign inter_9[388] = inter_8[388];
    assign inter_9[389] = inter_8[389];
    assign inter_9[390] = inter_8[390];
    assign inter_9[391] = inter_8[391];
    assign inter_9[392] = inter_8[392];
    assign inter_9[393] = inter_8[393];
    assign inter_9[394] = inter_8[394];
    assign inter_9[395] = inter_8[395];
    assign inter_9[396] = inter_8[396];
    assign inter_9[397] = inter_8[397];
    assign inter_9[398] = inter_8[398];
    assign inter_9[399] = inter_8[399];
    assign inter_9[400] = inter_8[400];
    assign inter_9[401] = inter_8[401];
    assign inter_9[402] = inter_8[402];
    assign inter_9[403] = inter_8[403];
    assign inter_9[404] = inter_8[404];
    assign inter_9[405] = inter_8[405];
    assign inter_9[406] = inter_8[406];
    assign inter_9[407] = inter_8[407];
    assign inter_9[408] = inter_8[408];
    assign inter_9[409] = inter_8[409];
    assign inter_9[410] = inter_8[410];
    assign inter_9[411] = inter_8[411];
    assign inter_9[412] = inter_8[412];
    assign inter_9[413] = inter_8[413];
    assign inter_9[414] = inter_8[414];
    assign inter_9[415] = inter_8[415];
    assign inter_9[416] = inter_8[416];
    assign inter_9[417] = inter_8[417];
    assign inter_9[418] = inter_8[418];
    assign inter_9[419] = inter_8[419];
    assign inter_9[420] = inter_8[420];
    assign inter_9[421] = inter_8[421];
    assign inter_9[422] = inter_8[422];
    assign inter_9[423] = inter_8[423];
    assign inter_9[424] = inter_8[424];
    assign inter_9[425] = inter_8[425];
    assign inter_9[426] = inter_8[426];
    assign inter_9[427] = inter_8[427];
    assign inter_9[428] = inter_8[428];
    assign inter_9[429] = inter_8[429];
    assign inter_9[430] = inter_8[430];
    assign inter_9[431] = inter_8[431];
    assign inter_9[432] = inter_8[432];
    assign inter_9[433] = inter_8[433];
    assign inter_9[434] = inter_8[434];
    assign inter_9[435] = inter_8[435];
    assign inter_9[436] = inter_8[436];
    assign inter_9[437] = inter_8[437];
    assign inter_9[438] = inter_8[438];
    assign inter_9[439] = inter_8[439];
    assign inter_9[440] = inter_8[440];
    assign inter_9[441] = inter_8[441];
    assign inter_9[442] = inter_8[442];
    assign inter_9[443] = inter_8[443];
    assign inter_9[444] = inter_8[444];
    assign inter_9[445] = inter_8[445];
    assign inter_9[446] = inter_8[446];
    assign inter_9[447] = inter_8[447];
    assign inter_9[448] = inter_8[448];
    assign inter_9[449] = inter_8[449];
    assign inter_9[450] = inter_8[450];
    assign inter_9[451] = inter_8[451];
    assign inter_9[452] = inter_8[452];
    assign inter_9[453] = inter_8[453];
    assign inter_9[454] = inter_8[454];
    assign inter_9[455] = inter_8[455];
    assign inter_9[456] = inter_8[456];
    assign inter_9[457] = inter_8[457];
    assign inter_9[458] = inter_8[458];
    assign inter_9[459] = inter_8[459];
    assign inter_9[460] = inter_8[460];
    assign inter_9[461] = inter_8[461];
    assign inter_9[462] = inter_8[462];
    assign inter_9[463] = inter_8[463];
    assign inter_9[464] = inter_8[464];
    assign inter_9[465] = inter_8[465];
    assign inter_9[466] = inter_8[466];
    assign inter_9[467] = inter_8[467];
    assign inter_9[468] = inter_8[468];
    assign inter_9[469] = inter_8[469];
    assign inter_9[470] = inter_8[470];
    assign inter_9[471] = inter_8[471];
    assign inter_9[472] = inter_8[472];
    assign inter_9[473] = inter_8[473];
    assign inter_9[474] = inter_8[474];
    assign inter_9[475] = inter_8[475];
    assign inter_9[476] = inter_8[476];
    assign inter_9[477] = inter_8[477];
    assign inter_9[478] = inter_8[478];
    assign inter_9[479] = inter_8[479];
    assign inter_9[480] = inter_8[480];
    assign inter_9[481] = inter_8[481];
    assign inter_9[482] = inter_8[482];
    assign inter_9[483] = inter_8[483];
    assign inter_9[484] = inter_8[484];
    assign inter_9[485] = inter_8[485];
    assign inter_9[486] = inter_8[486];
    assign inter_9[487] = inter_8[487];
    assign inter_9[488] = inter_8[488];
    assign inter_9[489] = inter_8[489];
    assign inter_9[490] = inter_8[490];
    assign inter_9[491] = inter_8[491];
    assign inter_9[492] = inter_8[492];
    assign inter_9[493] = inter_8[493];
    assign inter_9[494] = inter_8[494];
    assign inter_9[495] = inter_8[495];
    assign inter_9[496] = inter_8[496];
    assign inter_9[497] = inter_8[497];
    assign inter_9[498] = inter_8[498];
    assign inter_9[499] = inter_8[499];
    assign inter_9[500] = inter_8[500];
    assign inter_9[501] = inter_8[501];
    assign inter_9[502] = inter_8[502];
    assign inter_9[503] = inter_8[503];
    assign inter_9[504] = inter_8[504];
    assign inter_9[505] = inter_8[505];
    assign inter_9[506] = inter_8[506];
    assign inter_9[507] = inter_8[507];
    assign inter_9[508] = inter_8[508];
    assign inter_9[509] = inter_8[509];
    assign inter_9[510] = inter_8[510];
    assign inter_9[511] = inter_8[511];
    assign inter_9[512] = inter_8[512]^inter_8[768];
    assign inter_9[513] = inter_8[513]^inter_8[769];
    assign inter_9[514] = inter_8[514]^inter_8[770];
    assign inter_9[515] = inter_8[515]^inter_8[771];
    assign inter_9[516] = inter_8[516]^inter_8[772];
    assign inter_9[517] = inter_8[517]^inter_8[773];
    assign inter_9[518] = inter_8[518]^inter_8[774];
    assign inter_9[519] = inter_8[519]^inter_8[775];
    assign inter_9[520] = inter_8[520]^inter_8[776];
    assign inter_9[521] = inter_8[521]^inter_8[777];
    assign inter_9[522] = inter_8[522]^inter_8[778];
    assign inter_9[523] = inter_8[523]^inter_8[779];
    assign inter_9[524] = inter_8[524]^inter_8[780];
    assign inter_9[525] = inter_8[525]^inter_8[781];
    assign inter_9[526] = inter_8[526]^inter_8[782];
    assign inter_9[527] = inter_8[527]^inter_8[783];
    assign inter_9[528] = inter_8[528]^inter_8[784];
    assign inter_9[529] = inter_8[529]^inter_8[785];
    assign inter_9[530] = inter_8[530]^inter_8[786];
    assign inter_9[531] = inter_8[531]^inter_8[787];
    assign inter_9[532] = inter_8[532]^inter_8[788];
    assign inter_9[533] = inter_8[533]^inter_8[789];
    assign inter_9[534] = inter_8[534]^inter_8[790];
    assign inter_9[535] = inter_8[535]^inter_8[791];
    assign inter_9[536] = inter_8[536]^inter_8[792];
    assign inter_9[537] = inter_8[537]^inter_8[793];
    assign inter_9[538] = inter_8[538]^inter_8[794];
    assign inter_9[539] = inter_8[539]^inter_8[795];
    assign inter_9[540] = inter_8[540]^inter_8[796];
    assign inter_9[541] = inter_8[541]^inter_8[797];
    assign inter_9[542] = inter_8[542]^inter_8[798];
    assign inter_9[543] = inter_8[543]^inter_8[799];
    assign inter_9[544] = inter_8[544]^inter_8[800];
    assign inter_9[545] = inter_8[545]^inter_8[801];
    assign inter_9[546] = inter_8[546]^inter_8[802];
    assign inter_9[547] = inter_8[547]^inter_8[803];
    assign inter_9[548] = inter_8[548]^inter_8[804];
    assign inter_9[549] = inter_8[549]^inter_8[805];
    assign inter_9[550] = inter_8[550]^inter_8[806];
    assign inter_9[551] = inter_8[551]^inter_8[807];
    assign inter_9[552] = inter_8[552]^inter_8[808];
    assign inter_9[553] = inter_8[553]^inter_8[809];
    assign inter_9[554] = inter_8[554]^inter_8[810];
    assign inter_9[555] = inter_8[555]^inter_8[811];
    assign inter_9[556] = inter_8[556]^inter_8[812];
    assign inter_9[557] = inter_8[557]^inter_8[813];
    assign inter_9[558] = inter_8[558]^inter_8[814];
    assign inter_9[559] = inter_8[559]^inter_8[815];
    assign inter_9[560] = inter_8[560]^inter_8[816];
    assign inter_9[561] = inter_8[561]^inter_8[817];
    assign inter_9[562] = inter_8[562]^inter_8[818];
    assign inter_9[563] = inter_8[563]^inter_8[819];
    assign inter_9[564] = inter_8[564]^inter_8[820];
    assign inter_9[565] = inter_8[565]^inter_8[821];
    assign inter_9[566] = inter_8[566]^inter_8[822];
    assign inter_9[567] = inter_8[567]^inter_8[823];
    assign inter_9[568] = inter_8[568]^inter_8[824];
    assign inter_9[569] = inter_8[569]^inter_8[825];
    assign inter_9[570] = inter_8[570]^inter_8[826];
    assign inter_9[571] = inter_8[571]^inter_8[827];
    assign inter_9[572] = inter_8[572]^inter_8[828];
    assign inter_9[573] = inter_8[573]^inter_8[829];
    assign inter_9[574] = inter_8[574]^inter_8[830];
    assign inter_9[575] = inter_8[575]^inter_8[831];
    assign inter_9[576] = inter_8[576]^inter_8[832];
    assign inter_9[577] = inter_8[577]^inter_8[833];
    assign inter_9[578] = inter_8[578]^inter_8[834];
    assign inter_9[579] = inter_8[579]^inter_8[835];
    assign inter_9[580] = inter_8[580]^inter_8[836];
    assign inter_9[581] = inter_8[581]^inter_8[837];
    assign inter_9[582] = inter_8[582]^inter_8[838];
    assign inter_9[583] = inter_8[583]^inter_8[839];
    assign inter_9[584] = inter_8[584]^inter_8[840];
    assign inter_9[585] = inter_8[585]^inter_8[841];
    assign inter_9[586] = inter_8[586]^inter_8[842];
    assign inter_9[587] = inter_8[587]^inter_8[843];
    assign inter_9[588] = inter_8[588]^inter_8[844];
    assign inter_9[589] = inter_8[589]^inter_8[845];
    assign inter_9[590] = inter_8[590]^inter_8[846];
    assign inter_9[591] = inter_8[591]^inter_8[847];
    assign inter_9[592] = inter_8[592]^inter_8[848];
    assign inter_9[593] = inter_8[593]^inter_8[849];
    assign inter_9[594] = inter_8[594]^inter_8[850];
    assign inter_9[595] = inter_8[595]^inter_8[851];
    assign inter_9[596] = inter_8[596]^inter_8[852];
    assign inter_9[597] = inter_8[597]^inter_8[853];
    assign inter_9[598] = inter_8[598]^inter_8[854];
    assign inter_9[599] = inter_8[599]^inter_8[855];
    assign inter_9[600] = inter_8[600]^inter_8[856];
    assign inter_9[601] = inter_8[601]^inter_8[857];
    assign inter_9[602] = inter_8[602]^inter_8[858];
    assign inter_9[603] = inter_8[603]^inter_8[859];
    assign inter_9[604] = inter_8[604]^inter_8[860];
    assign inter_9[605] = inter_8[605]^inter_8[861];
    assign inter_9[606] = inter_8[606]^inter_8[862];
    assign inter_9[607] = inter_8[607]^inter_8[863];
    assign inter_9[608] = inter_8[608]^inter_8[864];
    assign inter_9[609] = inter_8[609]^inter_8[865];
    assign inter_9[610] = inter_8[610]^inter_8[866];
    assign inter_9[611] = inter_8[611]^inter_8[867];
    assign inter_9[612] = inter_8[612]^inter_8[868];
    assign inter_9[613] = inter_8[613]^inter_8[869];
    assign inter_9[614] = inter_8[614]^inter_8[870];
    assign inter_9[615] = inter_8[615]^inter_8[871];
    assign inter_9[616] = inter_8[616]^inter_8[872];
    assign inter_9[617] = inter_8[617]^inter_8[873];
    assign inter_9[618] = inter_8[618]^inter_8[874];
    assign inter_9[619] = inter_8[619]^inter_8[875];
    assign inter_9[620] = inter_8[620]^inter_8[876];
    assign inter_9[621] = inter_8[621]^inter_8[877];
    assign inter_9[622] = inter_8[622]^inter_8[878];
    assign inter_9[623] = inter_8[623]^inter_8[879];
    assign inter_9[624] = inter_8[624]^inter_8[880];
    assign inter_9[625] = inter_8[625]^inter_8[881];
    assign inter_9[626] = inter_8[626]^inter_8[882];
    assign inter_9[627] = inter_8[627]^inter_8[883];
    assign inter_9[628] = inter_8[628]^inter_8[884];
    assign inter_9[629] = inter_8[629]^inter_8[885];
    assign inter_9[630] = inter_8[630]^inter_8[886];
    assign inter_9[631] = inter_8[631]^inter_8[887];
    assign inter_9[632] = inter_8[632]^inter_8[888];
    assign inter_9[633] = inter_8[633]^inter_8[889];
    assign inter_9[634] = inter_8[634]^inter_8[890];
    assign inter_9[635] = inter_8[635]^inter_8[891];
    assign inter_9[636] = inter_8[636]^inter_8[892];
    assign inter_9[637] = inter_8[637]^inter_8[893];
    assign inter_9[638] = inter_8[638]^inter_8[894];
    assign inter_9[639] = inter_8[639]^inter_8[895];
    assign inter_9[640] = inter_8[640]^inter_8[896];
    assign inter_9[641] = inter_8[641]^inter_8[897];
    assign inter_9[642] = inter_8[642]^inter_8[898];
    assign inter_9[643] = inter_8[643]^inter_8[899];
    assign inter_9[644] = inter_8[644]^inter_8[900];
    assign inter_9[645] = inter_8[645]^inter_8[901];
    assign inter_9[646] = inter_8[646]^inter_8[902];
    assign inter_9[647] = inter_8[647]^inter_8[903];
    assign inter_9[648] = inter_8[648]^inter_8[904];
    assign inter_9[649] = inter_8[649]^inter_8[905];
    assign inter_9[650] = inter_8[650]^inter_8[906];
    assign inter_9[651] = inter_8[651]^inter_8[907];
    assign inter_9[652] = inter_8[652]^inter_8[908];
    assign inter_9[653] = inter_8[653]^inter_8[909];
    assign inter_9[654] = inter_8[654]^inter_8[910];
    assign inter_9[655] = inter_8[655]^inter_8[911];
    assign inter_9[656] = inter_8[656]^inter_8[912];
    assign inter_9[657] = inter_8[657]^inter_8[913];
    assign inter_9[658] = inter_8[658]^inter_8[914];
    assign inter_9[659] = inter_8[659]^inter_8[915];
    assign inter_9[660] = inter_8[660]^inter_8[916];
    assign inter_9[661] = inter_8[661]^inter_8[917];
    assign inter_9[662] = inter_8[662]^inter_8[918];
    assign inter_9[663] = inter_8[663]^inter_8[919];
    assign inter_9[664] = inter_8[664]^inter_8[920];
    assign inter_9[665] = inter_8[665]^inter_8[921];
    assign inter_9[666] = inter_8[666]^inter_8[922];
    assign inter_9[667] = inter_8[667]^inter_8[923];
    assign inter_9[668] = inter_8[668]^inter_8[924];
    assign inter_9[669] = inter_8[669]^inter_8[925];
    assign inter_9[670] = inter_8[670]^inter_8[926];
    assign inter_9[671] = inter_8[671]^inter_8[927];
    assign inter_9[672] = inter_8[672]^inter_8[928];
    assign inter_9[673] = inter_8[673]^inter_8[929];
    assign inter_9[674] = inter_8[674]^inter_8[930];
    assign inter_9[675] = inter_8[675]^inter_8[931];
    assign inter_9[676] = inter_8[676]^inter_8[932];
    assign inter_9[677] = inter_8[677]^inter_8[933];
    assign inter_9[678] = inter_8[678]^inter_8[934];
    assign inter_9[679] = inter_8[679]^inter_8[935];
    assign inter_9[680] = inter_8[680]^inter_8[936];
    assign inter_9[681] = inter_8[681]^inter_8[937];
    assign inter_9[682] = inter_8[682]^inter_8[938];
    assign inter_9[683] = inter_8[683]^inter_8[939];
    assign inter_9[684] = inter_8[684]^inter_8[940];
    assign inter_9[685] = inter_8[685]^inter_8[941];
    assign inter_9[686] = inter_8[686]^inter_8[942];
    assign inter_9[687] = inter_8[687]^inter_8[943];
    assign inter_9[688] = inter_8[688]^inter_8[944];
    assign inter_9[689] = inter_8[689]^inter_8[945];
    assign inter_9[690] = inter_8[690]^inter_8[946];
    assign inter_9[691] = inter_8[691]^inter_8[947];
    assign inter_9[692] = inter_8[692]^inter_8[948];
    assign inter_9[693] = inter_8[693]^inter_8[949];
    assign inter_9[694] = inter_8[694]^inter_8[950];
    assign inter_9[695] = inter_8[695]^inter_8[951];
    assign inter_9[696] = inter_8[696]^inter_8[952];
    assign inter_9[697] = inter_8[697]^inter_8[953];
    assign inter_9[698] = inter_8[698]^inter_8[954];
    assign inter_9[699] = inter_8[699]^inter_8[955];
    assign inter_9[700] = inter_8[700]^inter_8[956];
    assign inter_9[701] = inter_8[701]^inter_8[957];
    assign inter_9[702] = inter_8[702]^inter_8[958];
    assign inter_9[703] = inter_8[703]^inter_8[959];
    assign inter_9[704] = inter_8[704]^inter_8[960];
    assign inter_9[705] = inter_8[705]^inter_8[961];
    assign inter_9[706] = inter_8[706]^inter_8[962];
    assign inter_9[707] = inter_8[707]^inter_8[963];
    assign inter_9[708] = inter_8[708]^inter_8[964];
    assign inter_9[709] = inter_8[709]^inter_8[965];
    assign inter_9[710] = inter_8[710]^inter_8[966];
    assign inter_9[711] = inter_8[711]^inter_8[967];
    assign inter_9[712] = inter_8[712]^inter_8[968];
    assign inter_9[713] = inter_8[713]^inter_8[969];
    assign inter_9[714] = inter_8[714]^inter_8[970];
    assign inter_9[715] = inter_8[715]^inter_8[971];
    assign inter_9[716] = inter_8[716]^inter_8[972];
    assign inter_9[717] = inter_8[717]^inter_8[973];
    assign inter_9[718] = inter_8[718]^inter_8[974];
    assign inter_9[719] = inter_8[719]^inter_8[975];
    assign inter_9[720] = inter_8[720]^inter_8[976];
    assign inter_9[721] = inter_8[721]^inter_8[977];
    assign inter_9[722] = inter_8[722]^inter_8[978];
    assign inter_9[723] = inter_8[723]^inter_8[979];
    assign inter_9[724] = inter_8[724]^inter_8[980];
    assign inter_9[725] = inter_8[725]^inter_8[981];
    assign inter_9[726] = inter_8[726]^inter_8[982];
    assign inter_9[727] = inter_8[727]^inter_8[983];
    assign inter_9[728] = inter_8[728]^inter_8[984];
    assign inter_9[729] = inter_8[729]^inter_8[985];
    assign inter_9[730] = inter_8[730]^inter_8[986];
    assign inter_9[731] = inter_8[731]^inter_8[987];
    assign inter_9[732] = inter_8[732]^inter_8[988];
    assign inter_9[733] = inter_8[733]^inter_8[989];
    assign inter_9[734] = inter_8[734]^inter_8[990];
    assign inter_9[735] = inter_8[735]^inter_8[991];
    assign inter_9[736] = inter_8[736]^inter_8[992];
    assign inter_9[737] = inter_8[737]^inter_8[993];
    assign inter_9[738] = inter_8[738]^inter_8[994];
    assign inter_9[739] = inter_8[739]^inter_8[995];
    assign inter_9[740] = inter_8[740]^inter_8[996];
    assign inter_9[741] = inter_8[741]^inter_8[997];
    assign inter_9[742] = inter_8[742]^inter_8[998];
    assign inter_9[743] = inter_8[743]^inter_8[999];
    assign inter_9[744] = inter_8[744]^inter_8[1000];
    assign inter_9[745] = inter_8[745]^inter_8[1001];
    assign inter_9[746] = inter_8[746]^inter_8[1002];
    assign inter_9[747] = inter_8[747]^inter_8[1003];
    assign inter_9[748] = inter_8[748]^inter_8[1004];
    assign inter_9[749] = inter_8[749]^inter_8[1005];
    assign inter_9[750] = inter_8[750]^inter_8[1006];
    assign inter_9[751] = inter_8[751]^inter_8[1007];
    assign inter_9[752] = inter_8[752]^inter_8[1008];
    assign inter_9[753] = inter_8[753]^inter_8[1009];
    assign inter_9[754] = inter_8[754]^inter_8[1010];
    assign inter_9[755] = inter_8[755]^inter_8[1011];
    assign inter_9[756] = inter_8[756]^inter_8[1012];
    assign inter_9[757] = inter_8[757]^inter_8[1013];
    assign inter_9[758] = inter_8[758]^inter_8[1014];
    assign inter_9[759] = inter_8[759]^inter_8[1015];
    assign inter_9[760] = inter_8[760]^inter_8[1016];
    assign inter_9[761] = inter_8[761]^inter_8[1017];
    assign inter_9[762] = inter_8[762]^inter_8[1018];
    assign inter_9[763] = inter_8[763]^inter_8[1019];
    assign inter_9[764] = inter_8[764]^inter_8[1020];
    assign inter_9[765] = inter_8[765]^inter_8[1021];
    assign inter_9[766] = inter_8[766]^inter_8[1022];
    assign inter_9[767] = inter_8[767]^inter_8[1023];
    assign inter_9[768] = inter_8[768];
    assign inter_9[769] = inter_8[769];
    assign inter_9[770] = inter_8[770];
    assign inter_9[771] = inter_8[771];
    assign inter_9[772] = inter_8[772];
    assign inter_9[773] = inter_8[773];
    assign inter_9[774] = inter_8[774];
    assign inter_9[775] = inter_8[775];
    assign inter_9[776] = inter_8[776];
    assign inter_9[777] = inter_8[777];
    assign inter_9[778] = inter_8[778];
    assign inter_9[779] = inter_8[779];
    assign inter_9[780] = inter_8[780];
    assign inter_9[781] = inter_8[781];
    assign inter_9[782] = inter_8[782];
    assign inter_9[783] = inter_8[783];
    assign inter_9[784] = inter_8[784];
    assign inter_9[785] = inter_8[785];
    assign inter_9[786] = inter_8[786];
    assign inter_9[787] = inter_8[787];
    assign inter_9[788] = inter_8[788];
    assign inter_9[789] = inter_8[789];
    assign inter_9[790] = inter_8[790];
    assign inter_9[791] = inter_8[791];
    assign inter_9[792] = inter_8[792];
    assign inter_9[793] = inter_8[793];
    assign inter_9[794] = inter_8[794];
    assign inter_9[795] = inter_8[795];
    assign inter_9[796] = inter_8[796];
    assign inter_9[797] = inter_8[797];
    assign inter_9[798] = inter_8[798];
    assign inter_9[799] = inter_8[799];
    assign inter_9[800] = inter_8[800];
    assign inter_9[801] = inter_8[801];
    assign inter_9[802] = inter_8[802];
    assign inter_9[803] = inter_8[803];
    assign inter_9[804] = inter_8[804];
    assign inter_9[805] = inter_8[805];
    assign inter_9[806] = inter_8[806];
    assign inter_9[807] = inter_8[807];
    assign inter_9[808] = inter_8[808];
    assign inter_9[809] = inter_8[809];
    assign inter_9[810] = inter_8[810];
    assign inter_9[811] = inter_8[811];
    assign inter_9[812] = inter_8[812];
    assign inter_9[813] = inter_8[813];
    assign inter_9[814] = inter_8[814];
    assign inter_9[815] = inter_8[815];
    assign inter_9[816] = inter_8[816];
    assign inter_9[817] = inter_8[817];
    assign inter_9[818] = inter_8[818];
    assign inter_9[819] = inter_8[819];
    assign inter_9[820] = inter_8[820];
    assign inter_9[821] = inter_8[821];
    assign inter_9[822] = inter_8[822];
    assign inter_9[823] = inter_8[823];
    assign inter_9[824] = inter_8[824];
    assign inter_9[825] = inter_8[825];
    assign inter_9[826] = inter_8[826];
    assign inter_9[827] = inter_8[827];
    assign inter_9[828] = inter_8[828];
    assign inter_9[829] = inter_8[829];
    assign inter_9[830] = inter_8[830];
    assign inter_9[831] = inter_8[831];
    assign inter_9[832] = inter_8[832];
    assign inter_9[833] = inter_8[833];
    assign inter_9[834] = inter_8[834];
    assign inter_9[835] = inter_8[835];
    assign inter_9[836] = inter_8[836];
    assign inter_9[837] = inter_8[837];
    assign inter_9[838] = inter_8[838];
    assign inter_9[839] = inter_8[839];
    assign inter_9[840] = inter_8[840];
    assign inter_9[841] = inter_8[841];
    assign inter_9[842] = inter_8[842];
    assign inter_9[843] = inter_8[843];
    assign inter_9[844] = inter_8[844];
    assign inter_9[845] = inter_8[845];
    assign inter_9[846] = inter_8[846];
    assign inter_9[847] = inter_8[847];
    assign inter_9[848] = inter_8[848];
    assign inter_9[849] = inter_8[849];
    assign inter_9[850] = inter_8[850];
    assign inter_9[851] = inter_8[851];
    assign inter_9[852] = inter_8[852];
    assign inter_9[853] = inter_8[853];
    assign inter_9[854] = inter_8[854];
    assign inter_9[855] = inter_8[855];
    assign inter_9[856] = inter_8[856];
    assign inter_9[857] = inter_8[857];
    assign inter_9[858] = inter_8[858];
    assign inter_9[859] = inter_8[859];
    assign inter_9[860] = inter_8[860];
    assign inter_9[861] = inter_8[861];
    assign inter_9[862] = inter_8[862];
    assign inter_9[863] = inter_8[863];
    assign inter_9[864] = inter_8[864];
    assign inter_9[865] = inter_8[865];
    assign inter_9[866] = inter_8[866];
    assign inter_9[867] = inter_8[867];
    assign inter_9[868] = inter_8[868];
    assign inter_9[869] = inter_8[869];
    assign inter_9[870] = inter_8[870];
    assign inter_9[871] = inter_8[871];
    assign inter_9[872] = inter_8[872];
    assign inter_9[873] = inter_8[873];
    assign inter_9[874] = inter_8[874];
    assign inter_9[875] = inter_8[875];
    assign inter_9[876] = inter_8[876];
    assign inter_9[877] = inter_8[877];
    assign inter_9[878] = inter_8[878];
    assign inter_9[879] = inter_8[879];
    assign inter_9[880] = inter_8[880];
    assign inter_9[881] = inter_8[881];
    assign inter_9[882] = inter_8[882];
    assign inter_9[883] = inter_8[883];
    assign inter_9[884] = inter_8[884];
    assign inter_9[885] = inter_8[885];
    assign inter_9[886] = inter_8[886];
    assign inter_9[887] = inter_8[887];
    assign inter_9[888] = inter_8[888];
    assign inter_9[889] = inter_8[889];
    assign inter_9[890] = inter_8[890];
    assign inter_9[891] = inter_8[891];
    assign inter_9[892] = inter_8[892];
    assign inter_9[893] = inter_8[893];
    assign inter_9[894] = inter_8[894];
    assign inter_9[895] = inter_8[895];
    assign inter_9[896] = inter_8[896];
    assign inter_9[897] = inter_8[897];
    assign inter_9[898] = inter_8[898];
    assign inter_9[899] = inter_8[899];
    assign inter_9[900] = inter_8[900];
    assign inter_9[901] = inter_8[901];
    assign inter_9[902] = inter_8[902];
    assign inter_9[903] = inter_8[903];
    assign inter_9[904] = inter_8[904];
    assign inter_9[905] = inter_8[905];
    assign inter_9[906] = inter_8[906];
    assign inter_9[907] = inter_8[907];
    assign inter_9[908] = inter_8[908];
    assign inter_9[909] = inter_8[909];
    assign inter_9[910] = inter_8[910];
    assign inter_9[911] = inter_8[911];
    assign inter_9[912] = inter_8[912];
    assign inter_9[913] = inter_8[913];
    assign inter_9[914] = inter_8[914];
    assign inter_9[915] = inter_8[915];
    assign inter_9[916] = inter_8[916];
    assign inter_9[917] = inter_8[917];
    assign inter_9[918] = inter_8[918];
    assign inter_9[919] = inter_8[919];
    assign inter_9[920] = inter_8[920];
    assign inter_9[921] = inter_8[921];
    assign inter_9[922] = inter_8[922];
    assign inter_9[923] = inter_8[923];
    assign inter_9[924] = inter_8[924];
    assign inter_9[925] = inter_8[925];
    assign inter_9[926] = inter_8[926];
    assign inter_9[927] = inter_8[927];
    assign inter_9[928] = inter_8[928];
    assign inter_9[929] = inter_8[929];
    assign inter_9[930] = inter_8[930];
    assign inter_9[931] = inter_8[931];
    assign inter_9[932] = inter_8[932];
    assign inter_9[933] = inter_8[933];
    assign inter_9[934] = inter_8[934];
    assign inter_9[935] = inter_8[935];
    assign inter_9[936] = inter_8[936];
    assign inter_9[937] = inter_8[937];
    assign inter_9[938] = inter_8[938];
    assign inter_9[939] = inter_8[939];
    assign inter_9[940] = inter_8[940];
    assign inter_9[941] = inter_8[941];
    assign inter_9[942] = inter_8[942];
    assign inter_9[943] = inter_8[943];
    assign inter_9[944] = inter_8[944];
    assign inter_9[945] = inter_8[945];
    assign inter_9[946] = inter_8[946];
    assign inter_9[947] = inter_8[947];
    assign inter_9[948] = inter_8[948];
    assign inter_9[949] = inter_8[949];
    assign inter_9[950] = inter_8[950];
    assign inter_9[951] = inter_8[951];
    assign inter_9[952] = inter_8[952];
    assign inter_9[953] = inter_8[953];
    assign inter_9[954] = inter_8[954];
    assign inter_9[955] = inter_8[955];
    assign inter_9[956] = inter_8[956];
    assign inter_9[957] = inter_8[957];
    assign inter_9[958] = inter_8[958];
    assign inter_9[959] = inter_8[959];
    assign inter_9[960] = inter_8[960];
    assign inter_9[961] = inter_8[961];
    assign inter_9[962] = inter_8[962];
    assign inter_9[963] = inter_8[963];
    assign inter_9[964] = inter_8[964];
    assign inter_9[965] = inter_8[965];
    assign inter_9[966] = inter_8[966];
    assign inter_9[967] = inter_8[967];
    assign inter_9[968] = inter_8[968];
    assign inter_9[969] = inter_8[969];
    assign inter_9[970] = inter_8[970];
    assign inter_9[971] = inter_8[971];
    assign inter_9[972] = inter_8[972];
    assign inter_9[973] = inter_8[973];
    assign inter_9[974] = inter_8[974];
    assign inter_9[975] = inter_8[975];
    assign inter_9[976] = inter_8[976];
    assign inter_9[977] = inter_8[977];
    assign inter_9[978] = inter_8[978];
    assign inter_9[979] = inter_8[979];
    assign inter_9[980] = inter_8[980];
    assign inter_9[981] = inter_8[981];
    assign inter_9[982] = inter_8[982];
    assign inter_9[983] = inter_8[983];
    assign inter_9[984] = inter_8[984];
    assign inter_9[985] = inter_8[985];
    assign inter_9[986] = inter_8[986];
    assign inter_9[987] = inter_8[987];
    assign inter_9[988] = inter_8[988];
    assign inter_9[989] = inter_8[989];
    assign inter_9[990] = inter_8[990];
    assign inter_9[991] = inter_8[991];
    assign inter_9[992] = inter_8[992];
    assign inter_9[993] = inter_8[993];
    assign inter_9[994] = inter_8[994];
    assign inter_9[995] = inter_8[995];
    assign inter_9[996] = inter_8[996];
    assign inter_9[997] = inter_8[997];
    assign inter_9[998] = inter_8[998];
    assign inter_9[999] = inter_8[999];
    assign inter_9[1000] = inter_8[1000];
    assign inter_9[1001] = inter_8[1001];
    assign inter_9[1002] = inter_8[1002];
    assign inter_9[1003] = inter_8[1003];
    assign inter_9[1004] = inter_8[1004];
    assign inter_9[1005] = inter_8[1005];
    assign inter_9[1006] = inter_8[1006];
    assign inter_9[1007] = inter_8[1007];
    assign inter_9[1008] = inter_8[1008];
    assign inter_9[1009] = inter_8[1009];
    assign inter_9[1010] = inter_8[1010];
    assign inter_9[1011] = inter_8[1011];
    assign inter_9[1012] = inter_8[1012];
    assign inter_9[1013] = inter_8[1013];
    assign inter_9[1014] = inter_8[1014];
    assign inter_9[1015] = inter_8[1015];
    assign inter_9[1016] = inter_8[1016];
    assign inter_9[1017] = inter_8[1017];
    assign inter_9[1018] = inter_8[1018];
    assign inter_9[1019] = inter_8[1019];
    assign inter_9[1020] = inter_8[1020];
    assign inter_9[1021] = inter_8[1021];
    assign inter_9[1022] = inter_8[1022];
    assign inter_9[1023] = inter_8[1023];
    /***************************/
    assign inter_10[0] = inter_9[0]^inter_9[512];
    assign inter_10[1] = inter_9[1]^inter_9[513];
    assign inter_10[2] = inter_9[2]^inter_9[514];
    assign inter_10[3] = inter_9[3]^inter_9[515];
    assign inter_10[4] = inter_9[4]^inter_9[516];
    assign inter_10[5] = inter_9[5]^inter_9[517];
    assign inter_10[6] = inter_9[6]^inter_9[518];
    assign inter_10[7] = inter_9[7]^inter_9[519];
    assign inter_10[8] = inter_9[8]^inter_9[520];
    assign inter_10[9] = inter_9[9]^inter_9[521];
    assign inter_10[10] = inter_9[10]^inter_9[522];
    assign inter_10[11] = inter_9[11]^inter_9[523];
    assign inter_10[12] = inter_9[12]^inter_9[524];
    assign inter_10[13] = inter_9[13]^inter_9[525];
    assign inter_10[14] = inter_9[14]^inter_9[526];
    assign inter_10[15] = inter_9[15]^inter_9[527];
    assign inter_10[16] = inter_9[16]^inter_9[528];
    assign inter_10[17] = inter_9[17]^inter_9[529];
    assign inter_10[18] = inter_9[18]^inter_9[530];
    assign inter_10[19] = inter_9[19]^inter_9[531];
    assign inter_10[20] = inter_9[20]^inter_9[532];
    assign inter_10[21] = inter_9[21]^inter_9[533];
    assign inter_10[22] = inter_9[22]^inter_9[534];
    assign inter_10[23] = inter_9[23]^inter_9[535];
    assign inter_10[24] = inter_9[24]^inter_9[536];
    assign inter_10[25] = inter_9[25]^inter_9[537];
    assign inter_10[26] = inter_9[26]^inter_9[538];
    assign inter_10[27] = inter_9[27]^inter_9[539];
    assign inter_10[28] = inter_9[28]^inter_9[540];
    assign inter_10[29] = inter_9[29]^inter_9[541];
    assign inter_10[30] = inter_9[30]^inter_9[542];
    assign inter_10[31] = inter_9[31]^inter_9[543];
    assign inter_10[32] = inter_9[32]^inter_9[544];
    assign inter_10[33] = inter_9[33]^inter_9[545];
    assign inter_10[34] = inter_9[34]^inter_9[546];
    assign inter_10[35] = inter_9[35]^inter_9[547];
    assign inter_10[36] = inter_9[36]^inter_9[548];
    assign inter_10[37] = inter_9[37]^inter_9[549];
    assign inter_10[38] = inter_9[38]^inter_9[550];
    assign inter_10[39] = inter_9[39]^inter_9[551];
    assign inter_10[40] = inter_9[40]^inter_9[552];
    assign inter_10[41] = inter_9[41]^inter_9[553];
    assign inter_10[42] = inter_9[42]^inter_9[554];
    assign inter_10[43] = inter_9[43]^inter_9[555];
    assign inter_10[44] = inter_9[44]^inter_9[556];
    assign inter_10[45] = inter_9[45]^inter_9[557];
    assign inter_10[46] = inter_9[46]^inter_9[558];
    assign inter_10[47] = inter_9[47]^inter_9[559];
    assign inter_10[48] = inter_9[48]^inter_9[560];
    assign inter_10[49] = inter_9[49]^inter_9[561];
    assign inter_10[50] = inter_9[50]^inter_9[562];
    assign inter_10[51] = inter_9[51]^inter_9[563];
    assign inter_10[52] = inter_9[52]^inter_9[564];
    assign inter_10[53] = inter_9[53]^inter_9[565];
    assign inter_10[54] = inter_9[54]^inter_9[566];
    assign inter_10[55] = inter_9[55]^inter_9[567];
    assign inter_10[56] = inter_9[56]^inter_9[568];
    assign inter_10[57] = inter_9[57]^inter_9[569];
    assign inter_10[58] = inter_9[58]^inter_9[570];
    assign inter_10[59] = inter_9[59]^inter_9[571];
    assign inter_10[60] = inter_9[60]^inter_9[572];
    assign inter_10[61] = inter_9[61]^inter_9[573];
    assign inter_10[62] = inter_9[62]^inter_9[574];
    assign inter_10[63] = inter_9[63]^inter_9[575];
    assign inter_10[64] = inter_9[64]^inter_9[576];
    assign inter_10[65] = inter_9[65]^inter_9[577];
    assign inter_10[66] = inter_9[66]^inter_9[578];
    assign inter_10[67] = inter_9[67]^inter_9[579];
    assign inter_10[68] = inter_9[68]^inter_9[580];
    assign inter_10[69] = inter_9[69]^inter_9[581];
    assign inter_10[70] = inter_9[70]^inter_9[582];
    assign inter_10[71] = inter_9[71]^inter_9[583];
    assign inter_10[72] = inter_9[72]^inter_9[584];
    assign inter_10[73] = inter_9[73]^inter_9[585];
    assign inter_10[74] = inter_9[74]^inter_9[586];
    assign inter_10[75] = inter_9[75]^inter_9[587];
    assign inter_10[76] = inter_9[76]^inter_9[588];
    assign inter_10[77] = inter_9[77]^inter_9[589];
    assign inter_10[78] = inter_9[78]^inter_9[590];
    assign inter_10[79] = inter_9[79]^inter_9[591];
    assign inter_10[80] = inter_9[80]^inter_9[592];
    assign inter_10[81] = inter_9[81]^inter_9[593];
    assign inter_10[82] = inter_9[82]^inter_9[594];
    assign inter_10[83] = inter_9[83]^inter_9[595];
    assign inter_10[84] = inter_9[84]^inter_9[596];
    assign inter_10[85] = inter_9[85]^inter_9[597];
    assign inter_10[86] = inter_9[86]^inter_9[598];
    assign inter_10[87] = inter_9[87]^inter_9[599];
    assign inter_10[88] = inter_9[88]^inter_9[600];
    assign inter_10[89] = inter_9[89]^inter_9[601];
    assign inter_10[90] = inter_9[90]^inter_9[602];
    assign inter_10[91] = inter_9[91]^inter_9[603];
    assign inter_10[92] = inter_9[92]^inter_9[604];
    assign inter_10[93] = inter_9[93]^inter_9[605];
    assign inter_10[94] = inter_9[94]^inter_9[606];
    assign inter_10[95] = inter_9[95]^inter_9[607];
    assign inter_10[96] = inter_9[96]^inter_9[608];
    assign inter_10[97] = inter_9[97]^inter_9[609];
    assign inter_10[98] = inter_9[98]^inter_9[610];
    assign inter_10[99] = inter_9[99]^inter_9[611];
    assign inter_10[100] = inter_9[100]^inter_9[612];
    assign inter_10[101] = inter_9[101]^inter_9[613];
    assign inter_10[102] = inter_9[102]^inter_9[614];
    assign inter_10[103] = inter_9[103]^inter_9[615];
    assign inter_10[104] = inter_9[104]^inter_9[616];
    assign inter_10[105] = inter_9[105]^inter_9[617];
    assign inter_10[106] = inter_9[106]^inter_9[618];
    assign inter_10[107] = inter_9[107]^inter_9[619];
    assign inter_10[108] = inter_9[108]^inter_9[620];
    assign inter_10[109] = inter_9[109]^inter_9[621];
    assign inter_10[110] = inter_9[110]^inter_9[622];
    assign inter_10[111] = inter_9[111]^inter_9[623];
    assign inter_10[112] = inter_9[112]^inter_9[624];
    assign inter_10[113] = inter_9[113]^inter_9[625];
    assign inter_10[114] = inter_9[114]^inter_9[626];
    assign inter_10[115] = inter_9[115]^inter_9[627];
    assign inter_10[116] = inter_9[116]^inter_9[628];
    assign inter_10[117] = inter_9[117]^inter_9[629];
    assign inter_10[118] = inter_9[118]^inter_9[630];
    assign inter_10[119] = inter_9[119]^inter_9[631];
    assign inter_10[120] = inter_9[120]^inter_9[632];
    assign inter_10[121] = inter_9[121]^inter_9[633];
    assign inter_10[122] = inter_9[122]^inter_9[634];
    assign inter_10[123] = inter_9[123]^inter_9[635];
    assign inter_10[124] = inter_9[124]^inter_9[636];
    assign inter_10[125] = inter_9[125]^inter_9[637];
    assign inter_10[126] = inter_9[126]^inter_9[638];
    assign inter_10[127] = inter_9[127]^inter_9[639];
    assign inter_10[128] = inter_9[128]^inter_9[640];
    assign inter_10[129] = inter_9[129]^inter_9[641];
    assign inter_10[130] = inter_9[130]^inter_9[642];
    assign inter_10[131] = inter_9[131]^inter_9[643];
    assign inter_10[132] = inter_9[132]^inter_9[644];
    assign inter_10[133] = inter_9[133]^inter_9[645];
    assign inter_10[134] = inter_9[134]^inter_9[646];
    assign inter_10[135] = inter_9[135]^inter_9[647];
    assign inter_10[136] = inter_9[136]^inter_9[648];
    assign inter_10[137] = inter_9[137]^inter_9[649];
    assign inter_10[138] = inter_9[138]^inter_9[650];
    assign inter_10[139] = inter_9[139]^inter_9[651];
    assign inter_10[140] = inter_9[140]^inter_9[652];
    assign inter_10[141] = inter_9[141]^inter_9[653];
    assign inter_10[142] = inter_9[142]^inter_9[654];
    assign inter_10[143] = inter_9[143]^inter_9[655];
    assign inter_10[144] = inter_9[144]^inter_9[656];
    assign inter_10[145] = inter_9[145]^inter_9[657];
    assign inter_10[146] = inter_9[146]^inter_9[658];
    assign inter_10[147] = inter_9[147]^inter_9[659];
    assign inter_10[148] = inter_9[148]^inter_9[660];
    assign inter_10[149] = inter_9[149]^inter_9[661];
    assign inter_10[150] = inter_9[150]^inter_9[662];
    assign inter_10[151] = inter_9[151]^inter_9[663];
    assign inter_10[152] = inter_9[152]^inter_9[664];
    assign inter_10[153] = inter_9[153]^inter_9[665];
    assign inter_10[154] = inter_9[154]^inter_9[666];
    assign inter_10[155] = inter_9[155]^inter_9[667];
    assign inter_10[156] = inter_9[156]^inter_9[668];
    assign inter_10[157] = inter_9[157]^inter_9[669];
    assign inter_10[158] = inter_9[158]^inter_9[670];
    assign inter_10[159] = inter_9[159]^inter_9[671];
    assign inter_10[160] = inter_9[160]^inter_9[672];
    assign inter_10[161] = inter_9[161]^inter_9[673];
    assign inter_10[162] = inter_9[162]^inter_9[674];
    assign inter_10[163] = inter_9[163]^inter_9[675];
    assign inter_10[164] = inter_9[164]^inter_9[676];
    assign inter_10[165] = inter_9[165]^inter_9[677];
    assign inter_10[166] = inter_9[166]^inter_9[678];
    assign inter_10[167] = inter_9[167]^inter_9[679];
    assign inter_10[168] = inter_9[168]^inter_9[680];
    assign inter_10[169] = inter_9[169]^inter_9[681];
    assign inter_10[170] = inter_9[170]^inter_9[682];
    assign inter_10[171] = inter_9[171]^inter_9[683];
    assign inter_10[172] = inter_9[172]^inter_9[684];
    assign inter_10[173] = inter_9[173]^inter_9[685];
    assign inter_10[174] = inter_9[174]^inter_9[686];
    assign inter_10[175] = inter_9[175]^inter_9[687];
    assign inter_10[176] = inter_9[176]^inter_9[688];
    assign inter_10[177] = inter_9[177]^inter_9[689];
    assign inter_10[178] = inter_9[178]^inter_9[690];
    assign inter_10[179] = inter_9[179]^inter_9[691];
    assign inter_10[180] = inter_9[180]^inter_9[692];
    assign inter_10[181] = inter_9[181]^inter_9[693];
    assign inter_10[182] = inter_9[182]^inter_9[694];
    assign inter_10[183] = inter_9[183]^inter_9[695];
    assign inter_10[184] = inter_9[184]^inter_9[696];
    assign inter_10[185] = inter_9[185]^inter_9[697];
    assign inter_10[186] = inter_9[186]^inter_9[698];
    assign inter_10[187] = inter_9[187]^inter_9[699];
    assign inter_10[188] = inter_9[188]^inter_9[700];
    assign inter_10[189] = inter_9[189]^inter_9[701];
    assign inter_10[190] = inter_9[190]^inter_9[702];
    assign inter_10[191] = inter_9[191]^inter_9[703];
    assign inter_10[192] = inter_9[192]^inter_9[704];
    assign inter_10[193] = inter_9[193]^inter_9[705];
    assign inter_10[194] = inter_9[194]^inter_9[706];
    assign inter_10[195] = inter_9[195]^inter_9[707];
    assign inter_10[196] = inter_9[196]^inter_9[708];
    assign inter_10[197] = inter_9[197]^inter_9[709];
    assign inter_10[198] = inter_9[198]^inter_9[710];
    assign inter_10[199] = inter_9[199]^inter_9[711];
    assign inter_10[200] = inter_9[200]^inter_9[712];
    assign inter_10[201] = inter_9[201]^inter_9[713];
    assign inter_10[202] = inter_9[202]^inter_9[714];
    assign inter_10[203] = inter_9[203]^inter_9[715];
    assign inter_10[204] = inter_9[204]^inter_9[716];
    assign inter_10[205] = inter_9[205]^inter_9[717];
    assign inter_10[206] = inter_9[206]^inter_9[718];
    assign inter_10[207] = inter_9[207]^inter_9[719];
    assign inter_10[208] = inter_9[208]^inter_9[720];
    assign inter_10[209] = inter_9[209]^inter_9[721];
    assign inter_10[210] = inter_9[210]^inter_9[722];
    assign inter_10[211] = inter_9[211]^inter_9[723];
    assign inter_10[212] = inter_9[212]^inter_9[724];
    assign inter_10[213] = inter_9[213]^inter_9[725];
    assign inter_10[214] = inter_9[214]^inter_9[726];
    assign inter_10[215] = inter_9[215]^inter_9[727];
    assign inter_10[216] = inter_9[216]^inter_9[728];
    assign inter_10[217] = inter_9[217]^inter_9[729];
    assign inter_10[218] = inter_9[218]^inter_9[730];
    assign inter_10[219] = inter_9[219]^inter_9[731];
    assign inter_10[220] = inter_9[220]^inter_9[732];
    assign inter_10[221] = inter_9[221]^inter_9[733];
    assign inter_10[222] = inter_9[222]^inter_9[734];
    assign inter_10[223] = inter_9[223]^inter_9[735];
    assign inter_10[224] = inter_9[224]^inter_9[736];
    assign inter_10[225] = inter_9[225]^inter_9[737];
    assign inter_10[226] = inter_9[226]^inter_9[738];
    assign inter_10[227] = inter_9[227]^inter_9[739];
    assign inter_10[228] = inter_9[228]^inter_9[740];
    assign inter_10[229] = inter_9[229]^inter_9[741];
    assign inter_10[230] = inter_9[230]^inter_9[742];
    assign inter_10[231] = inter_9[231]^inter_9[743];
    assign inter_10[232] = inter_9[232]^inter_9[744];
    assign inter_10[233] = inter_9[233]^inter_9[745];
    assign inter_10[234] = inter_9[234]^inter_9[746];
    assign inter_10[235] = inter_9[235]^inter_9[747];
    assign inter_10[236] = inter_9[236]^inter_9[748];
    assign inter_10[237] = inter_9[237]^inter_9[749];
    assign inter_10[238] = inter_9[238]^inter_9[750];
    assign inter_10[239] = inter_9[239]^inter_9[751];
    assign inter_10[240] = inter_9[240]^inter_9[752];
    assign inter_10[241] = inter_9[241]^inter_9[753];
    assign inter_10[242] = inter_9[242]^inter_9[754];
    assign inter_10[243] = inter_9[243]^inter_9[755];
    assign inter_10[244] = inter_9[244]^inter_9[756];
    assign inter_10[245] = inter_9[245]^inter_9[757];
    assign inter_10[246] = inter_9[246]^inter_9[758];
    assign inter_10[247] = inter_9[247]^inter_9[759];
    assign inter_10[248] = inter_9[248]^inter_9[760];
    assign inter_10[249] = inter_9[249]^inter_9[761];
    assign inter_10[250] = inter_9[250]^inter_9[762];
    assign inter_10[251] = inter_9[251]^inter_9[763];
    assign inter_10[252] = inter_9[252]^inter_9[764];
    assign inter_10[253] = inter_9[253]^inter_9[765];
    assign inter_10[254] = inter_9[254]^inter_9[766];
    assign inter_10[255] = inter_9[255]^inter_9[767];
    assign inter_10[256] = inter_9[256]^inter_9[768];
    assign inter_10[257] = inter_9[257]^inter_9[769];
    assign inter_10[258] = inter_9[258]^inter_9[770];
    assign inter_10[259] = inter_9[259]^inter_9[771];
    assign inter_10[260] = inter_9[260]^inter_9[772];
    assign inter_10[261] = inter_9[261]^inter_9[773];
    assign inter_10[262] = inter_9[262]^inter_9[774];
    assign inter_10[263] = inter_9[263]^inter_9[775];
    assign inter_10[264] = inter_9[264]^inter_9[776];
    assign inter_10[265] = inter_9[265]^inter_9[777];
    assign inter_10[266] = inter_9[266]^inter_9[778];
    assign inter_10[267] = inter_9[267]^inter_9[779];
    assign inter_10[268] = inter_9[268]^inter_9[780];
    assign inter_10[269] = inter_9[269]^inter_9[781];
    assign inter_10[270] = inter_9[270]^inter_9[782];
    assign inter_10[271] = inter_9[271]^inter_9[783];
    assign inter_10[272] = inter_9[272]^inter_9[784];
    assign inter_10[273] = inter_9[273]^inter_9[785];
    assign inter_10[274] = inter_9[274]^inter_9[786];
    assign inter_10[275] = inter_9[275]^inter_9[787];
    assign inter_10[276] = inter_9[276]^inter_9[788];
    assign inter_10[277] = inter_9[277]^inter_9[789];
    assign inter_10[278] = inter_9[278]^inter_9[790];
    assign inter_10[279] = inter_9[279]^inter_9[791];
    assign inter_10[280] = inter_9[280]^inter_9[792];
    assign inter_10[281] = inter_9[281]^inter_9[793];
    assign inter_10[282] = inter_9[282]^inter_9[794];
    assign inter_10[283] = inter_9[283]^inter_9[795];
    assign inter_10[284] = inter_9[284]^inter_9[796];
    assign inter_10[285] = inter_9[285]^inter_9[797];
    assign inter_10[286] = inter_9[286]^inter_9[798];
    assign inter_10[287] = inter_9[287]^inter_9[799];
    assign inter_10[288] = inter_9[288]^inter_9[800];
    assign inter_10[289] = inter_9[289]^inter_9[801];
    assign inter_10[290] = inter_9[290]^inter_9[802];
    assign inter_10[291] = inter_9[291]^inter_9[803];
    assign inter_10[292] = inter_9[292]^inter_9[804];
    assign inter_10[293] = inter_9[293]^inter_9[805];
    assign inter_10[294] = inter_9[294]^inter_9[806];
    assign inter_10[295] = inter_9[295]^inter_9[807];
    assign inter_10[296] = inter_9[296]^inter_9[808];
    assign inter_10[297] = inter_9[297]^inter_9[809];
    assign inter_10[298] = inter_9[298]^inter_9[810];
    assign inter_10[299] = inter_9[299]^inter_9[811];
    assign inter_10[300] = inter_9[300]^inter_9[812];
    assign inter_10[301] = inter_9[301]^inter_9[813];
    assign inter_10[302] = inter_9[302]^inter_9[814];
    assign inter_10[303] = inter_9[303]^inter_9[815];
    assign inter_10[304] = inter_9[304]^inter_9[816];
    assign inter_10[305] = inter_9[305]^inter_9[817];
    assign inter_10[306] = inter_9[306]^inter_9[818];
    assign inter_10[307] = inter_9[307]^inter_9[819];
    assign inter_10[308] = inter_9[308]^inter_9[820];
    assign inter_10[309] = inter_9[309]^inter_9[821];
    assign inter_10[310] = inter_9[310]^inter_9[822];
    assign inter_10[311] = inter_9[311]^inter_9[823];
    assign inter_10[312] = inter_9[312]^inter_9[824];
    assign inter_10[313] = inter_9[313]^inter_9[825];
    assign inter_10[314] = inter_9[314]^inter_9[826];
    assign inter_10[315] = inter_9[315]^inter_9[827];
    assign inter_10[316] = inter_9[316]^inter_9[828];
    assign inter_10[317] = inter_9[317]^inter_9[829];
    assign inter_10[318] = inter_9[318]^inter_9[830];
    assign inter_10[319] = inter_9[319]^inter_9[831];
    assign inter_10[320] = inter_9[320]^inter_9[832];
    assign inter_10[321] = inter_9[321]^inter_9[833];
    assign inter_10[322] = inter_9[322]^inter_9[834];
    assign inter_10[323] = inter_9[323]^inter_9[835];
    assign inter_10[324] = inter_9[324]^inter_9[836];
    assign inter_10[325] = inter_9[325]^inter_9[837];
    assign inter_10[326] = inter_9[326]^inter_9[838];
    assign inter_10[327] = inter_9[327]^inter_9[839];
    assign inter_10[328] = inter_9[328]^inter_9[840];
    assign inter_10[329] = inter_9[329]^inter_9[841];
    assign inter_10[330] = inter_9[330]^inter_9[842];
    assign inter_10[331] = inter_9[331]^inter_9[843];
    assign inter_10[332] = inter_9[332]^inter_9[844];
    assign inter_10[333] = inter_9[333]^inter_9[845];
    assign inter_10[334] = inter_9[334]^inter_9[846];
    assign inter_10[335] = inter_9[335]^inter_9[847];
    assign inter_10[336] = inter_9[336]^inter_9[848];
    assign inter_10[337] = inter_9[337]^inter_9[849];
    assign inter_10[338] = inter_9[338]^inter_9[850];
    assign inter_10[339] = inter_9[339]^inter_9[851];
    assign inter_10[340] = inter_9[340]^inter_9[852];
    assign inter_10[341] = inter_9[341]^inter_9[853];
    assign inter_10[342] = inter_9[342]^inter_9[854];
    assign inter_10[343] = inter_9[343]^inter_9[855];
    assign inter_10[344] = inter_9[344]^inter_9[856];
    assign inter_10[345] = inter_9[345]^inter_9[857];
    assign inter_10[346] = inter_9[346]^inter_9[858];
    assign inter_10[347] = inter_9[347]^inter_9[859];
    assign inter_10[348] = inter_9[348]^inter_9[860];
    assign inter_10[349] = inter_9[349]^inter_9[861];
    assign inter_10[350] = inter_9[350]^inter_9[862];
    assign inter_10[351] = inter_9[351]^inter_9[863];
    assign inter_10[352] = inter_9[352]^inter_9[864];
    assign inter_10[353] = inter_9[353]^inter_9[865];
    assign inter_10[354] = inter_9[354]^inter_9[866];
    assign inter_10[355] = inter_9[355]^inter_9[867];
    assign inter_10[356] = inter_9[356]^inter_9[868];
    assign inter_10[357] = inter_9[357]^inter_9[869];
    assign inter_10[358] = inter_9[358]^inter_9[870];
    assign inter_10[359] = inter_9[359]^inter_9[871];
    assign inter_10[360] = inter_9[360]^inter_9[872];
    assign inter_10[361] = inter_9[361]^inter_9[873];
    assign inter_10[362] = inter_9[362]^inter_9[874];
    assign inter_10[363] = inter_9[363]^inter_9[875];
    assign inter_10[364] = inter_9[364]^inter_9[876];
    assign inter_10[365] = inter_9[365]^inter_9[877];
    assign inter_10[366] = inter_9[366]^inter_9[878];
    assign inter_10[367] = inter_9[367]^inter_9[879];
    assign inter_10[368] = inter_9[368]^inter_9[880];
    assign inter_10[369] = inter_9[369]^inter_9[881];
    assign inter_10[370] = inter_9[370]^inter_9[882];
    assign inter_10[371] = inter_9[371]^inter_9[883];
    assign inter_10[372] = inter_9[372]^inter_9[884];
    assign inter_10[373] = inter_9[373]^inter_9[885];
    assign inter_10[374] = inter_9[374]^inter_9[886];
    assign inter_10[375] = inter_9[375]^inter_9[887];
    assign inter_10[376] = inter_9[376]^inter_9[888];
    assign inter_10[377] = inter_9[377]^inter_9[889];
    assign inter_10[378] = inter_9[378]^inter_9[890];
    assign inter_10[379] = inter_9[379]^inter_9[891];
    assign inter_10[380] = inter_9[380]^inter_9[892];
    assign inter_10[381] = inter_9[381]^inter_9[893];
    assign inter_10[382] = inter_9[382]^inter_9[894];
    assign inter_10[383] = inter_9[383]^inter_9[895];
    assign inter_10[384] = inter_9[384]^inter_9[896];
    assign inter_10[385] = inter_9[385]^inter_9[897];
    assign inter_10[386] = inter_9[386]^inter_9[898];
    assign inter_10[387] = inter_9[387]^inter_9[899];
    assign inter_10[388] = inter_9[388]^inter_9[900];
    assign inter_10[389] = inter_9[389]^inter_9[901];
    assign inter_10[390] = inter_9[390]^inter_9[902];
    assign inter_10[391] = inter_9[391]^inter_9[903];
    assign inter_10[392] = inter_9[392]^inter_9[904];
    assign inter_10[393] = inter_9[393]^inter_9[905];
    assign inter_10[394] = inter_9[394]^inter_9[906];
    assign inter_10[395] = inter_9[395]^inter_9[907];
    assign inter_10[396] = inter_9[396]^inter_9[908];
    assign inter_10[397] = inter_9[397]^inter_9[909];
    assign inter_10[398] = inter_9[398]^inter_9[910];
    assign inter_10[399] = inter_9[399]^inter_9[911];
    assign inter_10[400] = inter_9[400]^inter_9[912];
    assign inter_10[401] = inter_9[401]^inter_9[913];
    assign inter_10[402] = inter_9[402]^inter_9[914];
    assign inter_10[403] = inter_9[403]^inter_9[915];
    assign inter_10[404] = inter_9[404]^inter_9[916];
    assign inter_10[405] = inter_9[405]^inter_9[917];
    assign inter_10[406] = inter_9[406]^inter_9[918];
    assign inter_10[407] = inter_9[407]^inter_9[919];
    assign inter_10[408] = inter_9[408]^inter_9[920];
    assign inter_10[409] = inter_9[409]^inter_9[921];
    assign inter_10[410] = inter_9[410]^inter_9[922];
    assign inter_10[411] = inter_9[411]^inter_9[923];
    assign inter_10[412] = inter_9[412]^inter_9[924];
    assign inter_10[413] = inter_9[413]^inter_9[925];
    assign inter_10[414] = inter_9[414]^inter_9[926];
    assign inter_10[415] = inter_9[415]^inter_9[927];
    assign inter_10[416] = inter_9[416]^inter_9[928];
    assign inter_10[417] = inter_9[417]^inter_9[929];
    assign inter_10[418] = inter_9[418]^inter_9[930];
    assign inter_10[419] = inter_9[419]^inter_9[931];
    assign inter_10[420] = inter_9[420]^inter_9[932];
    assign inter_10[421] = inter_9[421]^inter_9[933];
    assign inter_10[422] = inter_9[422]^inter_9[934];
    assign inter_10[423] = inter_9[423]^inter_9[935];
    assign inter_10[424] = inter_9[424]^inter_9[936];
    assign inter_10[425] = inter_9[425]^inter_9[937];
    assign inter_10[426] = inter_9[426]^inter_9[938];
    assign inter_10[427] = inter_9[427]^inter_9[939];
    assign inter_10[428] = inter_9[428]^inter_9[940];
    assign inter_10[429] = inter_9[429]^inter_9[941];
    assign inter_10[430] = inter_9[430]^inter_9[942];
    assign inter_10[431] = inter_9[431]^inter_9[943];
    assign inter_10[432] = inter_9[432]^inter_9[944];
    assign inter_10[433] = inter_9[433]^inter_9[945];
    assign inter_10[434] = inter_9[434]^inter_9[946];
    assign inter_10[435] = inter_9[435]^inter_9[947];
    assign inter_10[436] = inter_9[436]^inter_9[948];
    assign inter_10[437] = inter_9[437]^inter_9[949];
    assign inter_10[438] = inter_9[438]^inter_9[950];
    assign inter_10[439] = inter_9[439]^inter_9[951];
    assign inter_10[440] = inter_9[440]^inter_9[952];
    assign inter_10[441] = inter_9[441]^inter_9[953];
    assign inter_10[442] = inter_9[442]^inter_9[954];
    assign inter_10[443] = inter_9[443]^inter_9[955];
    assign inter_10[444] = inter_9[444]^inter_9[956];
    assign inter_10[445] = inter_9[445]^inter_9[957];
    assign inter_10[446] = inter_9[446]^inter_9[958];
    assign inter_10[447] = inter_9[447]^inter_9[959];
    assign inter_10[448] = inter_9[448]^inter_9[960];
    assign inter_10[449] = inter_9[449]^inter_9[961];
    assign inter_10[450] = inter_9[450]^inter_9[962];
    assign inter_10[451] = inter_9[451]^inter_9[963];
    assign inter_10[452] = inter_9[452]^inter_9[964];
    assign inter_10[453] = inter_9[453]^inter_9[965];
    assign inter_10[454] = inter_9[454]^inter_9[966];
    assign inter_10[455] = inter_9[455]^inter_9[967];
    assign inter_10[456] = inter_9[456]^inter_9[968];
    assign inter_10[457] = inter_9[457]^inter_9[969];
    assign inter_10[458] = inter_9[458]^inter_9[970];
    assign inter_10[459] = inter_9[459]^inter_9[971];
    assign inter_10[460] = inter_9[460]^inter_9[972];
    assign inter_10[461] = inter_9[461]^inter_9[973];
    assign inter_10[462] = inter_9[462]^inter_9[974];
    assign inter_10[463] = inter_9[463]^inter_9[975];
    assign inter_10[464] = inter_9[464]^inter_9[976];
    assign inter_10[465] = inter_9[465]^inter_9[977];
    assign inter_10[466] = inter_9[466]^inter_9[978];
    assign inter_10[467] = inter_9[467]^inter_9[979];
    assign inter_10[468] = inter_9[468]^inter_9[980];
    assign inter_10[469] = inter_9[469]^inter_9[981];
    assign inter_10[470] = inter_9[470]^inter_9[982];
    assign inter_10[471] = inter_9[471]^inter_9[983];
    assign inter_10[472] = inter_9[472]^inter_9[984];
    assign inter_10[473] = inter_9[473]^inter_9[985];
    assign inter_10[474] = inter_9[474]^inter_9[986];
    assign inter_10[475] = inter_9[475]^inter_9[987];
    assign inter_10[476] = inter_9[476]^inter_9[988];
    assign inter_10[477] = inter_9[477]^inter_9[989];
    assign inter_10[478] = inter_9[478]^inter_9[990];
    assign inter_10[479] = inter_9[479]^inter_9[991];
    assign inter_10[480] = inter_9[480]^inter_9[992];
    assign inter_10[481] = inter_9[481]^inter_9[993];
    assign inter_10[482] = inter_9[482]^inter_9[994];
    assign inter_10[483] = inter_9[483]^inter_9[995];
    assign inter_10[484] = inter_9[484]^inter_9[996];
    assign inter_10[485] = inter_9[485]^inter_9[997];
    assign inter_10[486] = inter_9[486]^inter_9[998];
    assign inter_10[487] = inter_9[487]^inter_9[999];
    assign inter_10[488] = inter_9[488]^inter_9[1000];
    assign inter_10[489] = inter_9[489]^inter_9[1001];
    assign inter_10[490] = inter_9[490]^inter_9[1002];
    assign inter_10[491] = inter_9[491]^inter_9[1003];
    assign inter_10[492] = inter_9[492]^inter_9[1004];
    assign inter_10[493] = inter_9[493]^inter_9[1005];
    assign inter_10[494] = inter_9[494]^inter_9[1006];
    assign inter_10[495] = inter_9[495]^inter_9[1007];
    assign inter_10[496] = inter_9[496]^inter_9[1008];
    assign inter_10[497] = inter_9[497]^inter_9[1009];
    assign inter_10[498] = inter_9[498]^inter_9[1010];
    assign inter_10[499] = inter_9[499]^inter_9[1011];
    assign inter_10[500] = inter_9[500]^inter_9[1012];
    assign inter_10[501] = inter_9[501]^inter_9[1013];
    assign inter_10[502] = inter_9[502]^inter_9[1014];
    assign inter_10[503] = inter_9[503]^inter_9[1015];
    assign inter_10[504] = inter_9[504]^inter_9[1016];
    assign inter_10[505] = inter_9[505]^inter_9[1017];
    assign inter_10[506] = inter_9[506]^inter_9[1018];
    assign inter_10[507] = inter_9[507]^inter_9[1019];
    assign inter_10[508] = inter_9[508]^inter_9[1020];
    assign inter_10[509] = inter_9[509]^inter_9[1021];
    assign inter_10[510] = inter_9[510]^inter_9[1022];
    assign inter_10[511] = inter_9[511]^inter_9[1023];
    assign inter_10[512] = inter_9[512];
    assign inter_10[513] = inter_9[513];
    assign inter_10[514] = inter_9[514];
    assign inter_10[515] = inter_9[515];
    assign inter_10[516] = inter_9[516];
    assign inter_10[517] = inter_9[517];
    assign inter_10[518] = inter_9[518];
    assign inter_10[519] = inter_9[519];
    assign inter_10[520] = inter_9[520];
    assign inter_10[521] = inter_9[521];
    assign inter_10[522] = inter_9[522];
    assign inter_10[523] = inter_9[523];
    assign inter_10[524] = inter_9[524];
    assign inter_10[525] = inter_9[525];
    assign inter_10[526] = inter_9[526];
    assign inter_10[527] = inter_9[527];
    assign inter_10[528] = inter_9[528];
    assign inter_10[529] = inter_9[529];
    assign inter_10[530] = inter_9[530];
    assign inter_10[531] = inter_9[531];
    assign inter_10[532] = inter_9[532];
    assign inter_10[533] = inter_9[533];
    assign inter_10[534] = inter_9[534];
    assign inter_10[535] = inter_9[535];
    assign inter_10[536] = inter_9[536];
    assign inter_10[537] = inter_9[537];
    assign inter_10[538] = inter_9[538];
    assign inter_10[539] = inter_9[539];
    assign inter_10[540] = inter_9[540];
    assign inter_10[541] = inter_9[541];
    assign inter_10[542] = inter_9[542];
    assign inter_10[543] = inter_9[543];
    assign inter_10[544] = inter_9[544];
    assign inter_10[545] = inter_9[545];
    assign inter_10[546] = inter_9[546];
    assign inter_10[547] = inter_9[547];
    assign inter_10[548] = inter_9[548];
    assign inter_10[549] = inter_9[549];
    assign inter_10[550] = inter_9[550];
    assign inter_10[551] = inter_9[551];
    assign inter_10[552] = inter_9[552];
    assign inter_10[553] = inter_9[553];
    assign inter_10[554] = inter_9[554];
    assign inter_10[555] = inter_9[555];
    assign inter_10[556] = inter_9[556];
    assign inter_10[557] = inter_9[557];
    assign inter_10[558] = inter_9[558];
    assign inter_10[559] = inter_9[559];
    assign inter_10[560] = inter_9[560];
    assign inter_10[561] = inter_9[561];
    assign inter_10[562] = inter_9[562];
    assign inter_10[563] = inter_9[563];
    assign inter_10[564] = inter_9[564];
    assign inter_10[565] = inter_9[565];
    assign inter_10[566] = inter_9[566];
    assign inter_10[567] = inter_9[567];
    assign inter_10[568] = inter_9[568];
    assign inter_10[569] = inter_9[569];
    assign inter_10[570] = inter_9[570];
    assign inter_10[571] = inter_9[571];
    assign inter_10[572] = inter_9[572];
    assign inter_10[573] = inter_9[573];
    assign inter_10[574] = inter_9[574];
    assign inter_10[575] = inter_9[575];
    assign inter_10[576] = inter_9[576];
    assign inter_10[577] = inter_9[577];
    assign inter_10[578] = inter_9[578];
    assign inter_10[579] = inter_9[579];
    assign inter_10[580] = inter_9[580];
    assign inter_10[581] = inter_9[581];
    assign inter_10[582] = inter_9[582];
    assign inter_10[583] = inter_9[583];
    assign inter_10[584] = inter_9[584];
    assign inter_10[585] = inter_9[585];
    assign inter_10[586] = inter_9[586];
    assign inter_10[587] = inter_9[587];
    assign inter_10[588] = inter_9[588];
    assign inter_10[589] = inter_9[589];
    assign inter_10[590] = inter_9[590];
    assign inter_10[591] = inter_9[591];
    assign inter_10[592] = inter_9[592];
    assign inter_10[593] = inter_9[593];
    assign inter_10[594] = inter_9[594];
    assign inter_10[595] = inter_9[595];
    assign inter_10[596] = inter_9[596];
    assign inter_10[597] = inter_9[597];
    assign inter_10[598] = inter_9[598];
    assign inter_10[599] = inter_9[599];
    assign inter_10[600] = inter_9[600];
    assign inter_10[601] = inter_9[601];
    assign inter_10[602] = inter_9[602];
    assign inter_10[603] = inter_9[603];
    assign inter_10[604] = inter_9[604];
    assign inter_10[605] = inter_9[605];
    assign inter_10[606] = inter_9[606];
    assign inter_10[607] = inter_9[607];
    assign inter_10[608] = inter_9[608];
    assign inter_10[609] = inter_9[609];
    assign inter_10[610] = inter_9[610];
    assign inter_10[611] = inter_9[611];
    assign inter_10[612] = inter_9[612];
    assign inter_10[613] = inter_9[613];
    assign inter_10[614] = inter_9[614];
    assign inter_10[615] = inter_9[615];
    assign inter_10[616] = inter_9[616];
    assign inter_10[617] = inter_9[617];
    assign inter_10[618] = inter_9[618];
    assign inter_10[619] = inter_9[619];
    assign inter_10[620] = inter_9[620];
    assign inter_10[621] = inter_9[621];
    assign inter_10[622] = inter_9[622];
    assign inter_10[623] = inter_9[623];
    assign inter_10[624] = inter_9[624];
    assign inter_10[625] = inter_9[625];
    assign inter_10[626] = inter_9[626];
    assign inter_10[627] = inter_9[627];
    assign inter_10[628] = inter_9[628];
    assign inter_10[629] = inter_9[629];
    assign inter_10[630] = inter_9[630];
    assign inter_10[631] = inter_9[631];
    assign inter_10[632] = inter_9[632];
    assign inter_10[633] = inter_9[633];
    assign inter_10[634] = inter_9[634];
    assign inter_10[635] = inter_9[635];
    assign inter_10[636] = inter_9[636];
    assign inter_10[637] = inter_9[637];
    assign inter_10[638] = inter_9[638];
    assign inter_10[639] = inter_9[639];
    assign inter_10[640] = inter_9[640];
    assign inter_10[641] = inter_9[641];
    assign inter_10[642] = inter_9[642];
    assign inter_10[643] = inter_9[643];
    assign inter_10[644] = inter_9[644];
    assign inter_10[645] = inter_9[645];
    assign inter_10[646] = inter_9[646];
    assign inter_10[647] = inter_9[647];
    assign inter_10[648] = inter_9[648];
    assign inter_10[649] = inter_9[649];
    assign inter_10[650] = inter_9[650];
    assign inter_10[651] = inter_9[651];
    assign inter_10[652] = inter_9[652];
    assign inter_10[653] = inter_9[653];
    assign inter_10[654] = inter_9[654];
    assign inter_10[655] = inter_9[655];
    assign inter_10[656] = inter_9[656];
    assign inter_10[657] = inter_9[657];
    assign inter_10[658] = inter_9[658];
    assign inter_10[659] = inter_9[659];
    assign inter_10[660] = inter_9[660];
    assign inter_10[661] = inter_9[661];
    assign inter_10[662] = inter_9[662];
    assign inter_10[663] = inter_9[663];
    assign inter_10[664] = inter_9[664];
    assign inter_10[665] = inter_9[665];
    assign inter_10[666] = inter_9[666];
    assign inter_10[667] = inter_9[667];
    assign inter_10[668] = inter_9[668];
    assign inter_10[669] = inter_9[669];
    assign inter_10[670] = inter_9[670];
    assign inter_10[671] = inter_9[671];
    assign inter_10[672] = inter_9[672];
    assign inter_10[673] = inter_9[673];
    assign inter_10[674] = inter_9[674];
    assign inter_10[675] = inter_9[675];
    assign inter_10[676] = inter_9[676];
    assign inter_10[677] = inter_9[677];
    assign inter_10[678] = inter_9[678];
    assign inter_10[679] = inter_9[679];
    assign inter_10[680] = inter_9[680];
    assign inter_10[681] = inter_9[681];
    assign inter_10[682] = inter_9[682];
    assign inter_10[683] = inter_9[683];
    assign inter_10[684] = inter_9[684];
    assign inter_10[685] = inter_9[685];
    assign inter_10[686] = inter_9[686];
    assign inter_10[687] = inter_9[687];
    assign inter_10[688] = inter_9[688];
    assign inter_10[689] = inter_9[689];
    assign inter_10[690] = inter_9[690];
    assign inter_10[691] = inter_9[691];
    assign inter_10[692] = inter_9[692];
    assign inter_10[693] = inter_9[693];
    assign inter_10[694] = inter_9[694];
    assign inter_10[695] = inter_9[695];
    assign inter_10[696] = inter_9[696];
    assign inter_10[697] = inter_9[697];
    assign inter_10[698] = inter_9[698];
    assign inter_10[699] = inter_9[699];
    assign inter_10[700] = inter_9[700];
    assign inter_10[701] = inter_9[701];
    assign inter_10[702] = inter_9[702];
    assign inter_10[703] = inter_9[703];
    assign inter_10[704] = inter_9[704];
    assign inter_10[705] = inter_9[705];
    assign inter_10[706] = inter_9[706];
    assign inter_10[707] = inter_9[707];
    assign inter_10[708] = inter_9[708];
    assign inter_10[709] = inter_9[709];
    assign inter_10[710] = inter_9[710];
    assign inter_10[711] = inter_9[711];
    assign inter_10[712] = inter_9[712];
    assign inter_10[713] = inter_9[713];
    assign inter_10[714] = inter_9[714];
    assign inter_10[715] = inter_9[715];
    assign inter_10[716] = inter_9[716];
    assign inter_10[717] = inter_9[717];
    assign inter_10[718] = inter_9[718];
    assign inter_10[719] = inter_9[719];
    assign inter_10[720] = inter_9[720];
    assign inter_10[721] = inter_9[721];
    assign inter_10[722] = inter_9[722];
    assign inter_10[723] = inter_9[723];
    assign inter_10[724] = inter_9[724];
    assign inter_10[725] = inter_9[725];
    assign inter_10[726] = inter_9[726];
    assign inter_10[727] = inter_9[727];
    assign inter_10[728] = inter_9[728];
    assign inter_10[729] = inter_9[729];
    assign inter_10[730] = inter_9[730];
    assign inter_10[731] = inter_9[731];
    assign inter_10[732] = inter_9[732];
    assign inter_10[733] = inter_9[733];
    assign inter_10[734] = inter_9[734];
    assign inter_10[735] = inter_9[735];
    assign inter_10[736] = inter_9[736];
    assign inter_10[737] = inter_9[737];
    assign inter_10[738] = inter_9[738];
    assign inter_10[739] = inter_9[739];
    assign inter_10[740] = inter_9[740];
    assign inter_10[741] = inter_9[741];
    assign inter_10[742] = inter_9[742];
    assign inter_10[743] = inter_9[743];
    assign inter_10[744] = inter_9[744];
    assign inter_10[745] = inter_9[745];
    assign inter_10[746] = inter_9[746];
    assign inter_10[747] = inter_9[747];
    assign inter_10[748] = inter_9[748];
    assign inter_10[749] = inter_9[749];
    assign inter_10[750] = inter_9[750];
    assign inter_10[751] = inter_9[751];
    assign inter_10[752] = inter_9[752];
    assign inter_10[753] = inter_9[753];
    assign inter_10[754] = inter_9[754];
    assign inter_10[755] = inter_9[755];
    assign inter_10[756] = inter_9[756];
    assign inter_10[757] = inter_9[757];
    assign inter_10[758] = inter_9[758];
    assign inter_10[759] = inter_9[759];
    assign inter_10[760] = inter_9[760];
    assign inter_10[761] = inter_9[761];
    assign inter_10[762] = inter_9[762];
    assign inter_10[763] = inter_9[763];
    assign inter_10[764] = inter_9[764];
    assign inter_10[765] = inter_9[765];
    assign inter_10[766] = inter_9[766];
    assign inter_10[767] = inter_9[767];
    assign inter_10[768] = inter_9[768];
    assign inter_10[769] = inter_9[769];
    assign inter_10[770] = inter_9[770];
    assign inter_10[771] = inter_9[771];
    assign inter_10[772] = inter_9[772];
    assign inter_10[773] = inter_9[773];
    assign inter_10[774] = inter_9[774];
    assign inter_10[775] = inter_9[775];
    assign inter_10[776] = inter_9[776];
    assign inter_10[777] = inter_9[777];
    assign inter_10[778] = inter_9[778];
    assign inter_10[779] = inter_9[779];
    assign inter_10[780] = inter_9[780];
    assign inter_10[781] = inter_9[781];
    assign inter_10[782] = inter_9[782];
    assign inter_10[783] = inter_9[783];
    assign inter_10[784] = inter_9[784];
    assign inter_10[785] = inter_9[785];
    assign inter_10[786] = inter_9[786];
    assign inter_10[787] = inter_9[787];
    assign inter_10[788] = inter_9[788];
    assign inter_10[789] = inter_9[789];
    assign inter_10[790] = inter_9[790];
    assign inter_10[791] = inter_9[791];
    assign inter_10[792] = inter_9[792];
    assign inter_10[793] = inter_9[793];
    assign inter_10[794] = inter_9[794];
    assign inter_10[795] = inter_9[795];
    assign inter_10[796] = inter_9[796];
    assign inter_10[797] = inter_9[797];
    assign inter_10[798] = inter_9[798];
    assign inter_10[799] = inter_9[799];
    assign inter_10[800] = inter_9[800];
    assign inter_10[801] = inter_9[801];
    assign inter_10[802] = inter_9[802];
    assign inter_10[803] = inter_9[803];
    assign inter_10[804] = inter_9[804];
    assign inter_10[805] = inter_9[805];
    assign inter_10[806] = inter_9[806];
    assign inter_10[807] = inter_9[807];
    assign inter_10[808] = inter_9[808];
    assign inter_10[809] = inter_9[809];
    assign inter_10[810] = inter_9[810];
    assign inter_10[811] = inter_9[811];
    assign inter_10[812] = inter_9[812];
    assign inter_10[813] = inter_9[813];
    assign inter_10[814] = inter_9[814];
    assign inter_10[815] = inter_9[815];
    assign inter_10[816] = inter_9[816];
    assign inter_10[817] = inter_9[817];
    assign inter_10[818] = inter_9[818];
    assign inter_10[819] = inter_9[819];
    assign inter_10[820] = inter_9[820];
    assign inter_10[821] = inter_9[821];
    assign inter_10[822] = inter_9[822];
    assign inter_10[823] = inter_9[823];
    assign inter_10[824] = inter_9[824];
    assign inter_10[825] = inter_9[825];
    assign inter_10[826] = inter_9[826];
    assign inter_10[827] = inter_9[827];
    assign inter_10[828] = inter_9[828];
    assign inter_10[829] = inter_9[829];
    assign inter_10[830] = inter_9[830];
    assign inter_10[831] = inter_9[831];
    assign inter_10[832] = inter_9[832];
    assign inter_10[833] = inter_9[833];
    assign inter_10[834] = inter_9[834];
    assign inter_10[835] = inter_9[835];
    assign inter_10[836] = inter_9[836];
    assign inter_10[837] = inter_9[837];
    assign inter_10[838] = inter_9[838];
    assign inter_10[839] = inter_9[839];
    assign inter_10[840] = inter_9[840];
    assign inter_10[841] = inter_9[841];
    assign inter_10[842] = inter_9[842];
    assign inter_10[843] = inter_9[843];
    assign inter_10[844] = inter_9[844];
    assign inter_10[845] = inter_9[845];
    assign inter_10[846] = inter_9[846];
    assign inter_10[847] = inter_9[847];
    assign inter_10[848] = inter_9[848];
    assign inter_10[849] = inter_9[849];
    assign inter_10[850] = inter_9[850];
    assign inter_10[851] = inter_9[851];
    assign inter_10[852] = inter_9[852];
    assign inter_10[853] = inter_9[853];
    assign inter_10[854] = inter_9[854];
    assign inter_10[855] = inter_9[855];
    assign inter_10[856] = inter_9[856];
    assign inter_10[857] = inter_9[857];
    assign inter_10[858] = inter_9[858];
    assign inter_10[859] = inter_9[859];
    assign inter_10[860] = inter_9[860];
    assign inter_10[861] = inter_9[861];
    assign inter_10[862] = inter_9[862];
    assign inter_10[863] = inter_9[863];
    assign inter_10[864] = inter_9[864];
    assign inter_10[865] = inter_9[865];
    assign inter_10[866] = inter_9[866];
    assign inter_10[867] = inter_9[867];
    assign inter_10[868] = inter_9[868];
    assign inter_10[869] = inter_9[869];
    assign inter_10[870] = inter_9[870];
    assign inter_10[871] = inter_9[871];
    assign inter_10[872] = inter_9[872];
    assign inter_10[873] = inter_9[873];
    assign inter_10[874] = inter_9[874];
    assign inter_10[875] = inter_9[875];
    assign inter_10[876] = inter_9[876];
    assign inter_10[877] = inter_9[877];
    assign inter_10[878] = inter_9[878];
    assign inter_10[879] = inter_9[879];
    assign inter_10[880] = inter_9[880];
    assign inter_10[881] = inter_9[881];
    assign inter_10[882] = inter_9[882];
    assign inter_10[883] = inter_9[883];
    assign inter_10[884] = inter_9[884];
    assign inter_10[885] = inter_9[885];
    assign inter_10[886] = inter_9[886];
    assign inter_10[887] = inter_9[887];
    assign inter_10[888] = inter_9[888];
    assign inter_10[889] = inter_9[889];
    assign inter_10[890] = inter_9[890];
    assign inter_10[891] = inter_9[891];
    assign inter_10[892] = inter_9[892];
    assign inter_10[893] = inter_9[893];
    assign inter_10[894] = inter_9[894];
    assign inter_10[895] = inter_9[895];
    assign inter_10[896] = inter_9[896];
    assign inter_10[897] = inter_9[897];
    assign inter_10[898] = inter_9[898];
    assign inter_10[899] = inter_9[899];
    assign inter_10[900] = inter_9[900];
    assign inter_10[901] = inter_9[901];
    assign inter_10[902] = inter_9[902];
    assign inter_10[903] = inter_9[903];
    assign inter_10[904] = inter_9[904];
    assign inter_10[905] = inter_9[905];
    assign inter_10[906] = inter_9[906];
    assign inter_10[907] = inter_9[907];
    assign inter_10[908] = inter_9[908];
    assign inter_10[909] = inter_9[909];
    assign inter_10[910] = inter_9[910];
    assign inter_10[911] = inter_9[911];
    assign inter_10[912] = inter_9[912];
    assign inter_10[913] = inter_9[913];
    assign inter_10[914] = inter_9[914];
    assign inter_10[915] = inter_9[915];
    assign inter_10[916] = inter_9[916];
    assign inter_10[917] = inter_9[917];
    assign inter_10[918] = inter_9[918];
    assign inter_10[919] = inter_9[919];
    assign inter_10[920] = inter_9[920];
    assign inter_10[921] = inter_9[921];
    assign inter_10[922] = inter_9[922];
    assign inter_10[923] = inter_9[923];
    assign inter_10[924] = inter_9[924];
    assign inter_10[925] = inter_9[925];
    assign inter_10[926] = inter_9[926];
    assign inter_10[927] = inter_9[927];
    assign inter_10[928] = inter_9[928];
    assign inter_10[929] = inter_9[929];
    assign inter_10[930] = inter_9[930];
    assign inter_10[931] = inter_9[931];
    assign inter_10[932] = inter_9[932];
    assign inter_10[933] = inter_9[933];
    assign inter_10[934] = inter_9[934];
    assign inter_10[935] = inter_9[935];
    assign inter_10[936] = inter_9[936];
    assign inter_10[937] = inter_9[937];
    assign inter_10[938] = inter_9[938];
    assign inter_10[939] = inter_9[939];
    assign inter_10[940] = inter_9[940];
    assign inter_10[941] = inter_9[941];
    assign inter_10[942] = inter_9[942];
    assign inter_10[943] = inter_9[943];
    assign inter_10[944] = inter_9[944];
    assign inter_10[945] = inter_9[945];
    assign inter_10[946] = inter_9[946];
    assign inter_10[947] = inter_9[947];
    assign inter_10[948] = inter_9[948];
    assign inter_10[949] = inter_9[949];
    assign inter_10[950] = inter_9[950];
    assign inter_10[951] = inter_9[951];
    assign inter_10[952] = inter_9[952];
    assign inter_10[953] = inter_9[953];
    assign inter_10[954] = inter_9[954];
    assign inter_10[955] = inter_9[955];
    assign inter_10[956] = inter_9[956];
    assign inter_10[957] = inter_9[957];
    assign inter_10[958] = inter_9[958];
    assign inter_10[959] = inter_9[959];
    assign inter_10[960] = inter_9[960];
    assign inter_10[961] = inter_9[961];
    assign inter_10[962] = inter_9[962];
    assign inter_10[963] = inter_9[963];
    assign inter_10[964] = inter_9[964];
    assign inter_10[965] = inter_9[965];
    assign inter_10[966] = inter_9[966];
    assign inter_10[967] = inter_9[967];
    assign inter_10[968] = inter_9[968];
    assign inter_10[969] = inter_9[969];
    assign inter_10[970] = inter_9[970];
    assign inter_10[971] = inter_9[971];
    assign inter_10[972] = inter_9[972];
    assign inter_10[973] = inter_9[973];
    assign inter_10[974] = inter_9[974];
    assign inter_10[975] = inter_9[975];
    assign inter_10[976] = inter_9[976];
    assign inter_10[977] = inter_9[977];
    assign inter_10[978] = inter_9[978];
    assign inter_10[979] = inter_9[979];
    assign inter_10[980] = inter_9[980];
    assign inter_10[981] = inter_9[981];
    assign inter_10[982] = inter_9[982];
    assign inter_10[983] = inter_9[983];
    assign inter_10[984] = inter_9[984];
    assign inter_10[985] = inter_9[985];
    assign inter_10[986] = inter_9[986];
    assign inter_10[987] = inter_9[987];
    assign inter_10[988] = inter_9[988];
    assign inter_10[989] = inter_9[989];
    assign inter_10[990] = inter_9[990];
    assign inter_10[991] = inter_9[991];
    assign inter_10[992] = inter_9[992];
    assign inter_10[993] = inter_9[993];
    assign inter_10[994] = inter_9[994];
    assign inter_10[995] = inter_9[995];
    assign inter_10[996] = inter_9[996];
    assign inter_10[997] = inter_9[997];
    assign inter_10[998] = inter_9[998];
    assign inter_10[999] = inter_9[999];
    assign inter_10[1000] = inter_9[1000];
    assign inter_10[1001] = inter_9[1001];
    assign inter_10[1002] = inter_9[1002];
    assign inter_10[1003] = inter_9[1003];
    assign inter_10[1004] = inter_9[1004];
    assign inter_10[1005] = inter_9[1005];
    assign inter_10[1006] = inter_9[1006];
    assign inter_10[1007] = inter_9[1007];
    assign inter_10[1008] = inter_9[1008];
    assign inter_10[1009] = inter_9[1009];
    assign inter_10[1010] = inter_9[1010];
    assign inter_10[1011] = inter_9[1011];
    assign inter_10[1012] = inter_9[1012];
    assign inter_10[1013] = inter_9[1013];
    assign inter_10[1014] = inter_9[1014];
    assign inter_10[1015] = inter_9[1015];
    assign inter_10[1016] = inter_9[1016];
    assign inter_10[1017] = inter_9[1017];
    assign inter_10[1018] = inter_9[1018];
    assign inter_10[1019] = inter_9[1019];
    assign inter_10[1020] = inter_9[1020];
    assign inter_10[1021] = inter_9[1021];
    assign inter_10[1022] = inter_9[1022];
    assign inter_10[1023] = inter_9[1023];
    /***************************/

  always @( posedge clk)
  begin
  if(rst)
  begin
   result = 0;
   end
   
  else 
  begin
  result = inter_10;
  end
  end
  piso ps(.clk(clk),.reset(reset),.parallel_in(result),.serial_out(result_s));
    
endmodule
